// Unpublished work. Copyright 2022 Siemens                         
// This material contains trade secrets or otherwise                
// confidential information owned by Siemens Industry Software Inc. 
// or its affiliates (collectively, "SISW"), or its licensors.      
// Access to and use of this information is strictly limited as     
// set forth in the Customer's applicable agreements with SISW.     
// This file was generated by profpga_brdgen version 14.0 
//   on Fri Dec 15 16:10:03 2023 

`timescale 1 ps / 1 ps

// Disable implicit declaration of wires
`default_nettype none

module top_fpga_mb1fb2
   (
    input  wire [7:0]  CLK_N,
    input  wire [7:0]  CLK_P,
    input  wire [7:0]  SYNC_N,
    input  wire [7:0]  SYNC_P,
    output wire [3:0]  SRC_CLK_N,
    output wire [3:0]  SRC_CLK_P,
    output wire [3:0]  SRC_SYNC_N,
    output wire [3:0]  SRC_SYNC_P,
    output wire [19:0] DMBI_F2H,
    input  wire [19:0] DMBI_H2F,
    input wire        mb1_FA2_TA0_CLKIO_N_0_mb1_FB2_TA2_CLKIO_N_7,
    input wire        mb1_FA2_TA0_CLKIO_N_1_mb1_FB2_TA2_CLKIO_N_6,
    input wire        mb1_FA2_TA0_CLKIO_N_2_mb1_FB2_TA2_CLKIO_N_4,
    input wire        mb1_FA2_TA0_CLKIO_N_3_mb1_FB2_TA2_CLKIO_N_3,
    input wire        mb1_FA2_TA0_CLKIO_N_4_mb1_FB2_TA2_CLKIO_N_2,
    input wire        mb1_FA2_TA0_CLKIO_N_5_mb1_FB2_TA2_IO_010,
    input wire        mb1_FA2_TA0_CLKIO_N_6_mb1_FB2_TA2_CLKIO_N_1,
    input wire        mb1_FA2_TA0_CLKIO_N_7_mb1_FB2_TA2_CLKIO_N_0,
    input wire        mb1_FA2_TA0_CLKIO_P_0_mb1_FB2_TA2_CLKIO_P_7,
    input wire        mb1_FA2_TA0_CLKIO_P_1_mb1_FB2_TA2_CLKIO_P_6,
    input wire        mb1_FA2_TA0_CLKIO_P_2_mb1_FB2_TA2_CLKIO_P_4,
    input wire        mb1_FA2_TA0_CLKIO_P_3_mb1_FB2_TA2_CLKIO_P_3,
    input wire        mb1_FA2_TA0_CLKIO_P_4_mb1_FB2_TA2_CLKIO_P_2,
    input wire        mb1_FA2_TA0_CLKIO_P_5_mb1_FB2_TA2_IO_011,
    input wire        mb1_FA2_TA0_CLKIO_P_6_mb1_FB2_TA2_CLKIO_P_1,
    input wire        mb1_FA2_TA0_CLKIO_P_7_mb1_FB2_TA2_CLKIO_P_0,
    input wire        mb1_FA2_TA0_IO_004_mb1_FB2_TA2_IO_006,
    input wire        mb1_FA2_TA0_IO_005_mb1_FB2_TA2_IO_007,
    input wire        mb1_FA2_TA0_IO_006_mb1_FB2_TA2_IO_004,
    input wire        mb1_FA2_TA0_IO_007_mb1_FB2_TA2_IO_005,
    input wire        mb1_FA2_TA0_IO_008_mb1_FB2_TA2_IO_022,
    input wire        mb1_FA2_TA0_IO_009_mb1_FB2_TA2_IO_023,
    input wire        mb1_FA2_TA0_IO_010_mb1_FB2_TA2_CLKIO_N_5,
    input wire        mb1_FA2_TA0_IO_011_mb1_FB2_TA2_CLKIO_P_5,
    input wire        mb1_FA2_TA0_IO_012_mb1_FB2_TA2_IO_012,
    input wire        mb1_FA2_TA0_IO_013_mb1_FB2_TA2_IO_013,
    input wire        mb1_FA2_TA0_IO_014_mb1_FB2_TA2_IO_016,
    input wire        mb1_FA2_TA0_IO_015_mb1_FB2_TA2_IO_017,
    input wire        mb1_FA2_TA0_IO_016_mb1_FB2_TA2_IO_014,
    input wire        mb1_FA2_TA0_IO_017_mb1_FB2_TA2_IO_015,
    input wire        mb1_FA2_TA0_IO_018_mb1_FB2_TA2_IO_032,
    input wire        mb1_FA2_TA0_IO_019_mb1_FB2_TA2_IO_033,
    input wire        mb1_FA2_TA0_IO_020_mb1_FB2_TA2_IO_030,
    input wire        mb1_FA2_TA0_IO_021_mb1_FB2_TA2_IO_031,
    input wire        mb1_FA2_TA0_IO_022_mb1_FB2_TA2_IO_008,
    input wire        mb1_FA2_TA0_IO_023_mb1_FB2_TA2_IO_009,
    input wire        mb1_FA2_TA0_IO_024_mb1_FB2_TA2_IO_026,
    input wire        mb1_FA2_TA0_IO_025_mb1_FB2_TA2_IO_027,
    input wire        mb1_FA2_TA0_IO_026_mb1_FB2_TA2_IO_024,
    input wire        mb1_FA2_TA0_IO_027_mb1_FB2_TA2_IO_025,
    input wire        mb1_FA2_TA0_IO_028_mb1_FB2_TA2_IO_042,
    input wire        mb1_FA2_TA0_IO_029_mb1_FB2_TA2_IO_043,
    input wire        mb1_FA2_TA0_IO_030_mb1_FB2_TA2_IO_020,
    input wire        mb1_FA2_TA0_IO_031_mb1_FB2_TA2_IO_021,
    input wire        mb1_FA2_TA0_IO_032_mb1_FB2_TA2_IO_018,
    input wire        mb1_FA2_TA0_IO_033_mb1_FB2_TA2_IO_019,
    input wire        mb1_FA2_TA0_IO_034_mb1_FB2_TA2_IO_036,
    input wire        mb1_FA2_TA0_IO_035_mb1_FB2_TA2_IO_037,
    input wire        mb1_FA2_TA0_IO_036_mb1_FB2_TA2_IO_034,
    input wire        mb1_FA2_TA0_IO_037_mb1_FB2_TA2_IO_035,
    input wire        mb1_FA2_TA0_IO_038_mb1_FB2_TA2_IO_052,
    input wire        mb1_FA2_TA0_IO_039_mb1_FB2_TA2_IO_053,
    input wire        mb1_FA2_TA0_IO_040_mb1_FB2_TA2_IO_050,
    input wire        mb1_FA2_TA0_IO_041_mb1_FB2_TA2_IO_051,
    input wire        mb1_FA2_TA0_IO_042_mb1_FB2_TA2_IO_028,
    input wire        mb1_FA2_TA0_IO_043_mb1_FB2_TA2_IO_029,
    input wire        mb1_FA2_TA0_IO_044_mb1_FB2_TA2_IO_046,
    input wire        mb1_FA2_TA0_IO_045_mb1_FB2_TA2_IO_047,
    input wire        mb1_FA2_TA0_IO_046_mb1_FB2_TA2_IO_044,
    input wire        mb1_FA2_TA0_IO_047_mb1_FB2_TA2_IO_045,
    input wire        mb1_FA2_TA0_IO_048_mb1_FB2_TA2_IO_062,
    input wire        mb1_FA2_TA0_IO_049_mb1_FB2_TA2_IO_063,
    input wire        mb1_FA2_TA0_IO_050_mb1_FB2_TA2_IO_040,
    input wire        mb1_FA2_TA0_IO_051_mb1_FB2_TA2_IO_041,
    input wire        mb1_FA2_TA0_IO_052_mb1_FB2_TA2_IO_038,
    input wire        mb1_FA2_TA0_IO_053_mb1_FB2_TA2_IO_039,
    input wire        mb1_FA2_TA0_IO_054_mb1_FB2_TA2_IO_056,
    input wire        mb1_FA2_TA0_IO_055_mb1_FB2_TA2_IO_057,
    input wire        mb1_FA2_TA0_IO_056_mb1_FB2_TA2_IO_054,
    input wire        mb1_FA2_TA0_IO_057_mb1_FB2_TA2_IO_055,
    input wire        mb1_FA2_TA0_IO_058_mb1_FB2_TA2_IO_072,
    input wire        mb1_FA2_TA0_IO_059_mb1_FB2_TA2_IO_073,
    input wire        mb1_FA2_TA0_IO_060_mb1_FB2_TA2_IO_070,
    input wire        mb1_FA2_TA0_IO_061_mb1_FB2_TA2_IO_071,
    input wire        mb1_FA2_TA0_IO_062_mb1_FB2_TA2_IO_048,
    input wire        mb1_FA2_TA0_IO_063_mb1_FB2_TA2_IO_049,
    input wire        mb1_FA2_TA0_IO_064_mb1_FB2_TA2_IO_066,
    input wire        mb1_FA2_TA0_IO_065_mb1_FB2_TA2_IO_067,
    input wire        mb1_FA2_TA0_IO_066_mb1_FB2_TA2_IO_064,
    input wire        mb1_FA2_TA0_IO_067_mb1_FB2_TA2_IO_065,
    input wire        mb1_FA2_TA0_IO_068_mb1_FB2_TA2_IO_082,
    input wire        mb1_FA2_TA0_IO_069_mb1_FB2_TA2_IO_083,
    input wire        mb1_FA2_TA0_IO_070_mb1_FB2_TA2_IO_060,
    input wire        mb1_FA2_TA0_IO_071_mb1_FB2_TA2_IO_061,
    input wire        mb1_FA2_TA0_IO_072_mb1_FB2_TA2_IO_058,
    input wire        mb1_FA2_TA0_IO_073_mb1_FB2_TA2_IO_059,
    input wire        mb1_FA2_TA0_IO_074_mb1_FB2_TA2_IO_076,
    input wire        mb1_FA2_TA0_IO_075_mb1_FB2_TA2_IO_077,
    input wire        mb1_FA2_TA0_IO_076_mb1_FB2_TA2_IO_074,
    input wire        mb1_FA2_TA0_IO_077_mb1_FB2_TA2_IO_075,
    input wire        mb1_FA2_TA0_IO_078_mb1_FB2_TA2_IO_092,
    input wire        mb1_FA2_TA0_IO_079_mb1_FB2_TA2_IO_093,
    input wire        mb1_FA2_TA0_IO_080_mb1_FB2_TA2_IO_090,
    input wire        mb1_FA2_TA0_IO_081_mb1_FB2_TA2_IO_091,
    input wire        mb1_FA2_TA0_IO_082_mb1_FB2_TA2_IO_068,
    input wire        mb1_FA2_TA0_IO_083_mb1_FB2_TA2_IO_069,
    input wire        mb1_FA2_TA0_IO_084_mb1_FB2_TA2_IO_086,
    input wire        mb1_FA2_TA0_IO_085_mb1_FB2_TA2_IO_087,
    input wire        mb1_FA2_TA0_IO_086_mb1_FB2_TA2_IO_084,
    input wire        mb1_FA2_TA0_IO_087_mb1_FB2_TA2_IO_085,
    input wire        mb1_FA2_TA0_IO_088_mb1_FB2_TA2_IO_102,
    input wire        mb1_FA2_TA0_IO_089_mb1_FB2_TA2_IO_103,
    input wire        mb1_FA2_TA0_IO_090_mb1_FB2_TA2_IO_080,
    input wire        mb1_FA2_TA0_IO_091_mb1_FB2_TA2_IO_081,
    input wire        mb1_FA2_TA0_IO_092_mb1_FB2_TA2_IO_078,
    input wire        mb1_FA2_TA0_IO_093_mb1_FB2_TA2_IO_079,
    input wire        mb1_FA2_TA0_IO_094_mb1_FB2_TA2_IO_096,
    input wire        mb1_FA2_TA0_IO_095_mb1_FB2_TA2_IO_097,
    input wire        mb1_FA2_TA0_IO_096_mb1_FB2_TA2_IO_094,
    input wire        mb1_FA2_TA0_IO_097_mb1_FB2_TA2_IO_095,
    input wire        mb1_FA2_TA0_IO_098_mb1_FB2_TA2_IO_112,
    input wire        mb1_FA2_TA0_IO_099_mb1_FB2_TA2_IO_113,
    input wire        mb1_FA2_TA0_IO_100_mb1_FB2_TA2_IO_110,
    input wire        mb1_FA2_TA0_IO_101_mb1_FB2_TA2_IO_111,
    input wire        mb1_FA2_TA0_IO_102_mb1_FB2_TA2_IO_088,
    input wire        mb1_FA2_TA0_IO_103_mb1_FB2_TA2_IO_089,
    input wire        mb1_FA2_TA0_IO_104_mb1_FB2_TA2_IO_106,
    input wire        mb1_FA2_TA0_IO_105_mb1_FB2_TA2_IO_107,
    input wire        mb1_FA2_TA0_IO_106_mb1_FB2_TA2_IO_104,
    input wire        mb1_FA2_TA0_IO_107_mb1_FB2_TA2_IO_105,
    input wire        mb1_FA2_TA0_IO_108_mb1_FB2_TA2_IO_122,
    input wire        mb1_FA2_TA0_IO_109_mb1_FB2_TA2_IO_123,
    input wire        mb1_FA2_TA0_IO_110_mb1_FB2_TA2_IO_100,
    input wire        mb1_FA2_TA0_IO_111_mb1_FB2_TA2_IO_101,
    input wire        mb1_FA2_TA0_IO_112_mb1_FB2_TA2_IO_098,
    input wire        mb1_FA2_TA0_IO_113_mb1_FB2_TA2_IO_099,
    input wire        mb1_FA2_TA0_IO_114_mb1_FB2_TA2_IO_116,
    input wire        mb1_FA2_TA0_IO_115_mb1_FB2_TA2_IO_117,
    input wire        mb1_FA2_TA0_IO_116_mb1_FB2_TA2_IO_114,
    input wire        mb1_FA2_TA0_IO_117_mb1_FB2_TA2_IO_115,
    input wire        mb1_FA2_TA0_IO_118_mb1_FB2_TA2_IO_132,
    input wire        mb1_FA2_TA0_IO_119_mb1_FB2_TA2_IO_133,
    input wire        mb1_FA2_TA0_IO_120_mb1_FB2_TA2_IO_130,
    input wire        mb1_FA2_TA0_IO_121_mb1_FB2_TA2_IO_131,
    input wire        mb1_FA2_TA0_IO_122_mb1_FB2_TA2_IO_108,
    input wire        mb1_FA2_TA0_IO_123_mb1_FB2_TA2_IO_109,
    input wire        mb1_FA2_TA0_IO_124_mb1_FB2_TA2_IO_126,
    input wire        mb1_FA2_TA0_IO_125_mb1_FB2_TA2_IO_127,
    input wire        mb1_FA2_TA0_IO_126_mb1_FB2_TA2_IO_124,
    input wire        mb1_FA2_TA0_IO_127_mb1_FB2_TA2_IO_125,
    input wire        mb1_FA2_TA0_IO_130_mb1_FB2_TA2_IO_120,
    input wire        mb1_FA2_TA0_IO_131_mb1_FB2_TA2_IO_121,
    input wire        mb1_FA2_TA0_IO_132_mb1_FB2_TA2_IO_118,
    input wire        mb1_FA2_TA0_IO_133_mb1_FB2_TA2_IO_119,
    input wire        mb1_FA2_TA0_IO_134_mb1_FB2_TA2_IO_136,
    input wire        mb1_FA2_TA0_IO_136_mb1_FB2_TA2_IO_134,
    input wire        mb1_FA2_BA0_CLKIO_N_0_mb1_FB2_TB0_CLKIO_N_7,
    input wire        mb1_FA2_BA0_CLKIO_N_1_mb1_FB2_TB0_CLKIO_N_6,
    input wire        mb1_FA2_BA0_CLKIO_N_2_mb1_FB2_TB0_CLKIO_N_4,
    input wire        mb1_FA2_BA0_CLKIO_N_3_mb1_FB2_TB0_CLKIO_N_3,
    input wire        mb1_FA2_BA0_CLKIO_N_4_mb1_FB2_TB0_CLKIO_N_2,
    input wire        mb1_FA2_BA0_CLKIO_N_5_mb1_FB2_TB0_IO_010,
    input wire        mb1_FA2_BA0_CLKIO_N_6_mb1_FB2_TB0_CLKIO_N_1,
    input wire        mb1_FA2_BA0_CLKIO_N_7_mb1_FB2_TB0_CLKIO_N_0,
    input wire        mb1_FA2_BA0_CLKIO_P_0_mb1_FB2_TB0_CLKIO_P_7,
    input wire        mb1_FA2_BA0_CLKIO_P_1_mb1_FB2_TB0_CLKIO_P_6,
    input wire        mb1_FA2_BA0_CLKIO_P_2_mb1_FB2_TB0_CLKIO_P_4,
    input wire        mb1_FA2_BA0_CLKIO_P_3_mb1_FB2_TB0_CLKIO_P_3,
    input wire        mb1_FA2_BA0_CLKIO_P_4_mb1_FB2_TB0_CLKIO_P_2,
    input wire        mb1_FA2_BA0_CLKIO_P_5_mb1_FB2_TB0_IO_011,
    input wire        mb1_FA2_BA0_CLKIO_P_6_mb1_FB2_TB0_CLKIO_P_1,
    input wire        mb1_FA2_BA0_CLKIO_P_7_mb1_FB2_TB0_CLKIO_P_0,
    input wire        mb1_FA2_BA0_IO_004_mb1_FB2_TB0_IO_006,
    input wire        mb1_FA2_BA0_IO_005_mb1_FB2_TB0_IO_007,
    input wire        mb1_FA2_BA0_IO_006_mb1_FB2_TB0_IO_004,
    input wire        mb1_FA2_BA0_IO_007_mb1_FB2_TB0_IO_005,
    input wire        mb1_FA2_BA0_IO_008_mb1_FB2_TB0_IO_022,
    input wire        mb1_FA2_BA0_IO_009_mb1_FB2_TB0_IO_023,
    input wire        mb1_FA2_BA0_IO_010_mb1_FB2_TB0_CLKIO_N_5,
    input wire        mb1_FA2_BA0_IO_011_mb1_FB2_TB0_CLKIO_P_5,
    input wire        mb1_FA2_BA0_IO_012_mb1_FB2_TB0_IO_012,
    input wire        mb1_FA2_BA0_IO_013_mb1_FB2_TB0_IO_013,
    input wire        mb1_FA2_BA0_IO_014_mb1_FB2_TB0_IO_016,
    input wire        mb1_FA2_BA0_IO_015_mb1_FB2_TB0_IO_017,
    input wire        mb1_FA2_BA0_IO_016_mb1_FB2_TB0_IO_014,
    input wire        mb1_FA2_BA0_IO_017_mb1_FB2_TB0_IO_015,
    input wire        mb1_FA2_BA0_IO_018_mb1_FB2_TB0_IO_032,
    input wire        mb1_FA2_BA0_IO_019_mb1_FB2_TB0_IO_033,
    input wire        mb1_FA2_BA0_IO_020_mb1_FB2_TB0_IO_030,
    input wire        mb1_FA2_BA0_IO_021_mb1_FB2_TB0_IO_031,
    input wire        mb1_FA2_BA0_IO_022_mb1_FB2_TB0_IO_008,
    input wire        mb1_FA2_BA0_IO_023_mb1_FB2_TB0_IO_009,
    input wire        mb1_FA2_BA0_IO_024_mb1_FB2_TB0_IO_026,
    input wire        mb1_FA2_BA0_IO_025_mb1_FB2_TB0_IO_027,
    input wire        mb1_FA2_BA0_IO_026_mb1_FB2_TB0_IO_024,
    input wire        mb1_FA2_BA0_IO_027_mb1_FB2_TB0_IO_025,
    input wire        mb1_FA2_BA0_IO_028_mb1_FB2_TB0_IO_042,
    input wire        mb1_FA2_BA0_IO_029_mb1_FB2_TB0_IO_043,
    input wire        mb1_FA2_BA0_IO_030_mb1_FB2_TB0_IO_020,
    input wire        mb1_FA2_BA0_IO_031_mb1_FB2_TB0_IO_021,
    input wire        mb1_FA2_BA0_IO_032_mb1_FB2_TB0_IO_018,
    input wire        mb1_FA2_BA0_IO_033_mb1_FB2_TB0_IO_019,
    input wire        mb1_FA2_BA0_IO_034_mb1_FB2_TB0_IO_036,
    input wire        mb1_FA2_BA0_IO_035_mb1_FB2_TB0_IO_037,
    input wire        mb1_FA2_BA0_IO_036_mb1_FB2_TB0_IO_034,
    input wire        mb1_FA2_BA0_IO_037_mb1_FB2_TB0_IO_035,
    input wire        mb1_FA2_BA0_IO_038_mb1_FB2_TB0_IO_052,
    input wire        mb1_FA2_BA0_IO_039_mb1_FB2_TB0_IO_053,
    input wire        mb1_FA2_BA0_IO_040_mb1_FB2_TB0_IO_050,
    input wire        mb1_FA2_BA0_IO_041_mb1_FB2_TB0_IO_051,
    input wire        mb1_FA2_BA0_IO_042_mb1_FB2_TB0_IO_028,
    input wire        mb1_FA2_BA0_IO_043_mb1_FB2_TB0_IO_029,
    input wire        mb1_FA2_BA0_IO_044_mb1_FB2_TB0_IO_046,
    input wire        mb1_FA2_BA0_IO_045_mb1_FB2_TB0_IO_047,
    input wire        mb1_FA2_BA0_IO_046_mb1_FB2_TB0_IO_044,
    input wire        mb1_FA2_BA0_IO_047_mb1_FB2_TB0_IO_045,
    input wire        mb1_FA2_BA0_IO_048_mb1_FB2_TB0_IO_062,
    input wire        mb1_FA2_BA0_IO_049_mb1_FB2_TB0_IO_063,
    input wire        mb1_FA2_BA0_IO_050_mb1_FB2_TB0_IO_040,
    input wire        mb1_FA2_BA0_IO_051_mb1_FB2_TB0_IO_041,
    input wire        mb1_FA2_BA0_IO_052_mb1_FB2_TB0_IO_038,
    input wire        mb1_FA2_BA0_IO_053_mb1_FB2_TB0_IO_039,
    input wire        mb1_FA2_BA0_IO_054_mb1_FB2_TB0_IO_056,
    input wire        mb1_FA2_BA0_IO_055_mb1_FB2_TB0_IO_057,
    input wire        mb1_FA2_BA0_IO_056_mb1_FB2_TB0_IO_054,
    input wire        mb1_FA2_BA0_IO_057_mb1_FB2_TB0_IO_055,
    input wire        mb1_FA2_BA0_IO_058_mb1_FB2_TB0_IO_072,
    input wire        mb1_FA2_BA0_IO_059_mb1_FB2_TB0_IO_073,
    input wire        mb1_FA2_BA0_IO_060_mb1_FB2_TB0_IO_070,
    input wire        mb1_FA2_BA0_IO_061_mb1_FB2_TB0_IO_071,
    input wire        mb1_FA2_BA0_IO_062_mb1_FB2_TB0_IO_048,
    input wire        mb1_FA2_BA0_IO_063_mb1_FB2_TB0_IO_049,
    input wire        mb1_FA2_BA0_IO_064_mb1_FB2_TB0_IO_066,
    input wire        mb1_FA2_BA0_IO_065_mb1_FB2_TB0_IO_067,
    input wire        mb1_FA2_BA0_IO_066_mb1_FB2_TB0_IO_064,
    input wire        mb1_FA2_BA0_IO_067_mb1_FB2_TB0_IO_065,
    input wire        mb1_FA2_BA0_IO_068_mb1_FB2_TB0_IO_082,
    input wire        mb1_FA2_BA0_IO_069_mb1_FB2_TB0_IO_083,
    input wire        mb1_FA2_BA0_IO_070_mb1_FB2_TB0_IO_060,
    input wire        mb1_FA2_BA0_IO_071_mb1_FB2_TB0_IO_061,
    input wire        mb1_FA2_BA0_IO_072_mb1_FB2_TB0_IO_058,
    input wire        mb1_FA2_BA0_IO_073_mb1_FB2_TB0_IO_059,
    input wire        mb1_FA2_BA0_IO_074_mb1_FB2_TB0_IO_076,
    input wire        mb1_FA2_BA0_IO_075_mb1_FB2_TB0_IO_077,
    input wire        mb1_FA2_BA0_IO_076_mb1_FB2_TB0_IO_074,
    input wire        mb1_FA2_BA0_IO_077_mb1_FB2_TB0_IO_075,
    input wire        mb1_FA2_BA0_IO_078_mb1_FB2_TB0_IO_092,
    input wire        mb1_FA2_BA0_IO_079_mb1_FB2_TB0_IO_093,
    input wire        mb1_FA2_BA0_IO_080_mb1_FB2_TB0_IO_090,
    input wire        mb1_FA2_BA0_IO_081_mb1_FB2_TB0_IO_091,
    input wire        mb1_FA2_BA0_IO_082_mb1_FB2_TB0_IO_068,
    input wire        mb1_FA2_BA0_IO_083_mb1_FB2_TB0_IO_069,
    input wire        mb1_FA2_BA0_IO_084_mb1_FB2_TB0_IO_086,
    input wire        mb1_FA2_BA0_IO_085_mb1_FB2_TB0_IO_087,
    input wire        mb1_FA2_BA0_IO_086_mb1_FB2_TB0_IO_084,
    input wire        mb1_FA2_BA0_IO_087_mb1_FB2_TB0_IO_085,
    input wire        mb1_FA2_BA0_IO_088_mb1_FB2_TB0_IO_102,
    input wire        mb1_FA2_BA0_IO_089_mb1_FB2_TB0_IO_103,
    input wire        mb1_FA2_BA0_IO_090_mb1_FB2_TB0_IO_080,
    input wire        mb1_FA2_BA0_IO_091_mb1_FB2_TB0_IO_081,
    input wire        mb1_FA2_BA0_IO_092_mb1_FB2_TB0_IO_078,
    input wire        mb1_FA2_BA0_IO_093_mb1_FB2_TB0_IO_079,
    input wire        mb1_FA2_BA0_IO_094_mb1_FB2_TB0_IO_096,
    input wire        mb1_FA2_BA0_IO_095_mb1_FB2_TB0_IO_097,
    input wire        mb1_FA2_BA0_IO_096_mb1_FB2_TB0_IO_094,
    input wire        mb1_FA2_BA0_IO_097_mb1_FB2_TB0_IO_095,
    input wire        mb1_FA2_BA0_IO_098_mb1_FB2_TB0_IO_112,
    input wire        mb1_FA2_BA0_IO_099_mb1_FB2_TB0_IO_113,
    input wire        mb1_FA2_BA0_IO_100_mb1_FB2_TB0_IO_110,
    input wire        mb1_FA2_BA0_IO_101_mb1_FB2_TB0_IO_111,
    input wire        mb1_FA2_BA0_IO_102_mb1_FB2_TB0_IO_088,
    input wire        mb1_FA2_BA0_IO_103_mb1_FB2_TB0_IO_089,
    input wire        mb1_FA2_BA0_IO_104_mb1_FB2_TB0_IO_106,
    input wire        mb1_FA2_BA0_IO_105_mb1_FB2_TB0_IO_107,
    input wire        mb1_FA2_BA0_IO_106_mb1_FB2_TB0_IO_104,
    input wire        mb1_FA2_BA0_IO_107_mb1_FB2_TB0_IO_105,
    input wire        mb1_FA2_BA0_IO_108_mb1_FB2_TB0_IO_122,
    input wire        mb1_FA2_BA0_IO_109_mb1_FB2_TB0_IO_123,
    input wire        mb1_FA2_BA0_IO_110_mb1_FB2_TB0_IO_100,
    input wire        mb1_FA2_BA0_IO_111_mb1_FB2_TB0_IO_101,
    input wire        mb1_FA2_BA0_IO_112_mb1_FB2_TB0_IO_098,
    input wire        mb1_FA2_BA0_IO_113_mb1_FB2_TB0_IO_099,
    input wire        mb1_FA2_BA0_IO_114_mb1_FB2_TB0_IO_116,
    input wire        mb1_FA2_BA0_IO_115_mb1_FB2_TB0_IO_117,
    input wire        mb1_FA2_BA0_IO_116_mb1_FB2_TB0_IO_114,
    input wire        mb1_FA2_BA0_IO_117_mb1_FB2_TB0_IO_115,
    input wire        mb1_FA2_BA0_IO_118_mb1_FB2_TB0_IO_132,
    input wire        mb1_FA2_BA0_IO_119_mb1_FB2_TB0_IO_133,
    input wire        mb1_FA2_BA0_IO_120_mb1_FB2_TB0_IO_130,
    input wire        mb1_FA2_BA0_IO_121_mb1_FB2_TB0_IO_131,
    input wire        mb1_FA2_BA0_IO_122_mb1_FB2_TB0_IO_108,
    input wire        mb1_FA2_BA0_IO_123_mb1_FB2_TB0_IO_109,
    input wire        mb1_FA2_BA0_IO_124_mb1_FB2_TB0_IO_126,
    input wire        mb1_FA2_BA0_IO_125_mb1_FB2_TB0_IO_127,
    input wire        mb1_FA2_BA0_IO_126_mb1_FB2_TB0_IO_124,
    input wire        mb1_FA2_BA0_IO_127_mb1_FB2_TB0_IO_125,
    input wire        mb1_FA2_BA0_IO_130_mb1_FB2_TB0_IO_120,
    input wire        mb1_FA2_BA0_IO_131_mb1_FB2_TB0_IO_121,
    input wire        mb1_FA2_BA0_IO_132_mb1_FB2_TB0_IO_118,
    input wire        mb1_FA2_BA0_IO_133_mb1_FB2_TB0_IO_119,
    input wire        mb1_FA2_BA0_IO_134_mb1_FB2_TB0_IO_136,
    input wire        mb1_FA2_BA0_IO_136_mb1_FB2_TB0_IO_134,
    input wire        mb1_FA2_TA2_CLKIO_N_0_mb1_FB2_TB1_CLKIO_N_7,
    input wire        mb1_FA2_TA2_CLKIO_N_1_mb1_FB2_TB1_CLKIO_N_6,
    input wire        mb1_FA2_TA2_CLKIO_N_2_mb1_FB2_TB1_CLKIO_N_4,
    input wire        mb1_FA2_TA2_CLKIO_N_3_mb1_FB2_TB1_CLKIO_N_3,
    input wire        mb1_FA2_TA2_CLKIO_N_4_mb1_FB2_TB1_CLKIO_N_2,
    input wire        mb1_FA2_TA2_CLKIO_N_5_mb1_FB2_TB1_IO_010,
    input wire        mb1_FA2_TA2_CLKIO_N_6_mb1_FB2_TB1_CLKIO_N_1,
    input wire        mb1_FA2_TA2_CLKIO_N_7_mb1_FB2_TB1_CLKIO_N_0,
    input wire        mb1_FA2_TA2_CLKIO_P_0_mb1_FB2_TB1_CLKIO_P_7,
    input wire        mb1_FA2_TA2_CLKIO_P_1_mb1_FB2_TB1_CLKIO_P_6,
    input wire        mb1_FA2_TA2_CLKIO_P_2_mb1_FB2_TB1_CLKIO_P_4,
    input wire        mb1_FA2_TA2_CLKIO_P_3_mb1_FB2_TB1_CLKIO_P_3,
    input wire        mb1_FA2_TA2_CLKIO_P_4_mb1_FB2_TB1_CLKIO_P_2,
    input wire        mb1_FA2_TA2_CLKIO_P_5_mb1_FB2_TB1_IO_011,
    input wire        mb1_FA2_TA2_CLKIO_P_6_mb1_FB2_TB1_CLKIO_P_1,
    input wire        mb1_FA2_TA2_CLKIO_P_7_mb1_FB2_TB1_CLKIO_P_0,
    input wire        mb1_FA2_TA2_IO_004_mb1_FB2_TB1_IO_006,
    input wire        mb1_FA2_TA2_IO_005_mb1_FB2_TB1_IO_007,
    input wire        mb1_FA2_TA2_IO_006_mb1_FB2_TB1_IO_004,
    input wire        mb1_FA2_TA2_IO_007_mb1_FB2_TB1_IO_005,
    input wire        mb1_FA2_TA2_IO_008_mb1_FB2_TB1_IO_022,
    input wire        mb1_FA2_TA2_IO_009_mb1_FB2_TB1_IO_023,
    input wire        mb1_FA2_TA2_IO_010_mb1_FB2_TB1_CLKIO_N_5,
    input wire        mb1_FA2_TA2_IO_011_mb1_FB2_TB1_CLKIO_P_5,
    input wire        mb1_FA2_TA2_IO_012_mb1_FB2_TB1_IO_012,
    input wire        mb1_FA2_TA2_IO_013_mb1_FB2_TB1_IO_013,
    input wire        mb1_FA2_TA2_IO_014_mb1_FB2_TB1_IO_016,
    input wire        mb1_FA2_TA2_IO_015_mb1_FB2_TB1_IO_017,
    input wire        mb1_FA2_TA2_IO_016_mb1_FB2_TB1_IO_014,
    input wire        mb1_FA2_TA2_IO_017_mb1_FB2_TB1_IO_015,
    input wire        mb1_FA2_TA2_IO_018_mb1_FB2_TB1_IO_032,
    input wire        mb1_FA2_TA2_IO_019_mb1_FB2_TB1_IO_033,
    input wire        mb1_FA2_TA2_IO_020_mb1_FB2_TB1_IO_030,
    input wire        mb1_FA2_TA2_IO_021_mb1_FB2_TB1_IO_031,
    input wire        mb1_FA2_TA2_IO_022_mb1_FB2_TB1_IO_008,
    input wire        mb1_FA2_TA2_IO_023_mb1_FB2_TB1_IO_009,
    input wire        mb1_FA2_TA2_IO_024_mb1_FB2_TB1_IO_026,
    input wire        mb1_FA2_TA2_IO_025_mb1_FB2_TB1_IO_027,
    input wire        mb1_FA2_TA2_IO_026_mb1_FB2_TB1_IO_024,
    input wire        mb1_FA2_TA2_IO_027_mb1_FB2_TB1_IO_025,
    input wire        mb1_FA2_TA2_IO_028_mb1_FB2_TB1_IO_042,
    input wire        mb1_FA2_TA2_IO_029_mb1_FB2_TB1_IO_043,
    input wire        mb1_FA2_TA2_IO_030_mb1_FB2_TB1_IO_020,
    input wire        mb1_FA2_TA2_IO_031_mb1_FB2_TB1_IO_021,
    input wire        mb1_FA2_TA2_IO_032_mb1_FB2_TB1_IO_018,
    input wire        mb1_FA2_TA2_IO_033_mb1_FB2_TB1_IO_019,
    input wire        mb1_FA2_TA2_IO_034_mb1_FB2_TB1_IO_036,
    input wire        mb1_FA2_TA2_IO_035_mb1_FB2_TB1_IO_037,
    input wire        mb1_FA2_TA2_IO_036_mb1_FB2_TB1_IO_034,
    input wire        mb1_FA2_TA2_IO_037_mb1_FB2_TB1_IO_035,
    input wire        mb1_FA2_TA2_IO_038_mb1_FB2_TB1_IO_052,
    input wire        mb1_FA2_TA2_IO_039_mb1_FB2_TB1_IO_053,
    input wire        mb1_FA2_TA2_IO_040_mb1_FB2_TB1_IO_050,
    input wire        mb1_FA2_TA2_IO_041_mb1_FB2_TB1_IO_051,
    input wire        mb1_FA2_TA2_IO_042_mb1_FB2_TB1_IO_028,
    input wire        mb1_FA2_TA2_IO_043_mb1_FB2_TB1_IO_029,
    input wire        mb1_FA2_TA2_IO_044_mb1_FB2_TB1_IO_046,
    input wire        mb1_FA2_TA2_IO_045_mb1_FB2_TB1_IO_047,
    input wire        mb1_FA2_TA2_IO_046_mb1_FB2_TB1_IO_044,
    input wire        mb1_FA2_TA2_IO_047_mb1_FB2_TB1_IO_045,
    input wire        mb1_FA2_TA2_IO_048_mb1_FB2_TB1_IO_062,
    input wire        mb1_FA2_TA2_IO_049_mb1_FB2_TB1_IO_063,
    input wire        mb1_FA2_TA2_IO_050_mb1_FB2_TB1_IO_040,
    input wire        mb1_FA2_TA2_IO_051_mb1_FB2_TB1_IO_041,
    input wire        mb1_FA2_TA2_IO_052_mb1_FB2_TB1_IO_038,
    input wire        mb1_FA2_TA2_IO_053_mb1_FB2_TB1_IO_039,
    input wire        mb1_FA2_TA2_IO_054_mb1_FB2_TB1_IO_056,
    input wire        mb1_FA2_TA2_IO_055_mb1_FB2_TB1_IO_057,
    input wire        mb1_FA2_TA2_IO_056_mb1_FB2_TB1_IO_054,
    input wire        mb1_FA2_TA2_IO_057_mb1_FB2_TB1_IO_055,
    input wire        mb1_FA2_TA2_IO_058_mb1_FB2_TB1_IO_072,
    input wire        mb1_FA2_TA2_IO_059_mb1_FB2_TB1_IO_073,
    input wire        mb1_FA2_TA2_IO_060_mb1_FB2_TB1_IO_070,
    input wire        mb1_FA2_TA2_IO_061_mb1_FB2_TB1_IO_071,
    input wire        mb1_FA2_TA2_IO_062_mb1_FB2_TB1_IO_048,
    input wire        mb1_FA2_TA2_IO_063_mb1_FB2_TB1_IO_049,
    input wire        mb1_FA2_TA2_IO_064_mb1_FB2_TB1_IO_066,
    input wire        mb1_FA2_TA2_IO_065_mb1_FB2_TB1_IO_067,
    input wire        mb1_FA2_TA2_IO_066_mb1_FB2_TB1_IO_064,
    input wire        mb1_FA2_TA2_IO_067_mb1_FB2_TB1_IO_065,
    input wire        mb1_FA2_TA2_IO_068_mb1_FB2_TB1_IO_082,
    input wire        mb1_FA2_TA2_IO_069_mb1_FB2_TB1_IO_083,
    input wire        mb1_FA2_TA2_IO_070_mb1_FB2_TB1_IO_060,
    input wire        mb1_FA2_TA2_IO_071_mb1_FB2_TB1_IO_061,
    input wire        mb1_FA2_TA2_IO_072_mb1_FB2_TB1_IO_058,
    input wire        mb1_FA2_TA2_IO_073_mb1_FB2_TB1_IO_059,
    input wire        mb1_FA2_TA2_IO_074_mb1_FB2_TB1_IO_076,
    input wire        mb1_FA2_TA2_IO_075_mb1_FB2_TB1_IO_077,
    input wire        mb1_FA2_TA2_IO_076_mb1_FB2_TB1_IO_074,
    input wire        mb1_FA2_TA2_IO_077_mb1_FB2_TB1_IO_075,
    input wire        mb1_FA2_TA2_IO_078_mb1_FB2_TB1_IO_092,
    input wire        mb1_FA2_TA2_IO_079_mb1_FB2_TB1_IO_093,
    input wire        mb1_FA2_TA2_IO_080_mb1_FB2_TB1_IO_090,
    input wire        mb1_FA2_TA2_IO_081_mb1_FB2_TB1_IO_091,
    input wire        mb1_FA2_TA2_IO_082_mb1_FB2_TB1_IO_068,
    input wire        mb1_FA2_TA2_IO_083_mb1_FB2_TB1_IO_069,
    input wire        mb1_FA2_TA2_IO_084_mb1_FB2_TB1_IO_086,
    input wire        mb1_FA2_TA2_IO_085_mb1_FB2_TB1_IO_087,
    input wire        mb1_FA2_TA2_IO_086_mb1_FB2_TB1_IO_084,
    input wire        mb1_FA2_TA2_IO_087_mb1_FB2_TB1_IO_085,
    input wire        mb1_FA2_TA2_IO_088_mb1_FB2_TB1_IO_102,
    input wire        mb1_FA2_TA2_IO_089_mb1_FB2_TB1_IO_103,
    input wire        mb1_FA2_TA2_IO_090_mb1_FB2_TB1_IO_080,
    input wire        mb1_FA2_TA2_IO_091_mb1_FB2_TB1_IO_081,
    input wire        mb1_FA2_TA2_IO_092_mb1_FB2_TB1_IO_078,
    input wire        mb1_FA2_TA2_IO_093_mb1_FB2_TB1_IO_079,
    input wire        mb1_FA2_TA2_IO_094_mb1_FB2_TB1_IO_096,
    input wire        mb1_FA2_TA2_IO_095_mb1_FB2_TB1_IO_097,
    input wire        mb1_FA2_TA2_IO_096_mb1_FB2_TB1_IO_094,
    input wire        mb1_FA2_TA2_IO_097_mb1_FB2_TB1_IO_095,
    input wire        mb1_FA2_TA2_IO_098_mb1_FB2_TB1_IO_112,
    input wire        mb1_FA2_TA2_IO_099_mb1_FB2_TB1_IO_113,
    input wire        mb1_FA2_TA2_IO_100_mb1_FB2_TB1_IO_110,
    input wire        mb1_FA2_TA2_IO_101_mb1_FB2_TB1_IO_111,
    input wire        mb1_FA2_TA2_IO_102_mb1_FB2_TB1_IO_088,
    input wire        mb1_FA2_TA2_IO_103_mb1_FB2_TB1_IO_089,
    input wire        mb1_FA2_TA2_IO_104_mb1_FB2_TB1_IO_106,
    input wire        mb1_FA2_TA2_IO_105_mb1_FB2_TB1_IO_107,
    input wire        mb1_FA2_TA2_IO_106_mb1_FB2_TB1_IO_104,
    input wire        mb1_FA2_TA2_IO_107_mb1_FB2_TB1_IO_105,
    input wire        mb1_FA2_TA2_IO_108_mb1_FB2_TB1_IO_122,
    input wire        mb1_FA2_TA2_IO_109_mb1_FB2_TB1_IO_123,
    input wire        mb1_FA2_TA2_IO_110_mb1_FB2_TB1_IO_100,
    input wire        mb1_FA2_TA2_IO_111_mb1_FB2_TB1_IO_101,
    input wire        mb1_FA2_TA2_IO_112_mb1_FB2_TB1_IO_098,
    input wire        mb1_FA2_TA2_IO_113_mb1_FB2_TB1_IO_099,
    input wire        mb1_FA2_TA2_IO_114_mb1_FB2_TB1_IO_116,
    input wire        mb1_FA2_TA2_IO_115_mb1_FB2_TB1_IO_117,
    input wire        mb1_FA2_TA2_IO_116_mb1_FB2_TB1_IO_114,
    input wire        mb1_FA2_TA2_IO_117_mb1_FB2_TB1_IO_115,
    input wire        mb1_FA2_TA2_IO_118_mb1_FB2_TB1_IO_132,
    input wire        mb1_FA2_TA2_IO_119_mb1_FB2_TB1_IO_133,
    input wire        mb1_FA2_TA2_IO_120_mb1_FB2_TB1_IO_130,
    input wire        mb1_FA2_TA2_IO_121_mb1_FB2_TB1_IO_131,
    input wire        mb1_FA2_TA2_IO_122_mb1_FB2_TB1_IO_108,
    input wire        mb1_FA2_TA2_IO_123_mb1_FB2_TB1_IO_109,
    input wire        mb1_FA2_TA2_IO_124_mb1_FB2_TB1_IO_126,
    input wire        mb1_FA2_TA2_IO_125_mb1_FB2_TB1_IO_127,
    input wire        mb1_FA2_TA2_IO_126_mb1_FB2_TB1_IO_124,
    input wire        mb1_FA2_TA2_IO_127_mb1_FB2_TB1_IO_125,
    input wire        mb1_FA2_TA2_IO_130_mb1_FB2_TB1_IO_120,
    input wire        mb1_FA2_TA2_IO_131_mb1_FB2_TB1_IO_121,
    input wire        mb1_FA2_TA2_IO_132_mb1_FB2_TB1_IO_118,
    input wire        mb1_FA2_TA2_IO_133_mb1_FB2_TB1_IO_119,
    input wire        mb1_FA2_TA2_IO_134_mb1_FB2_TB1_IO_136,
    input wire        mb1_FA2_TA2_IO_136_mb1_FB2_TB1_IO_134,
    input wire        mb1_FA2_TB2_CLKIO_N_0_mb1_FB2_TB2_CLKIO_N_7,
    input wire        mb1_FA2_TB2_CLKIO_N_1_mb1_FB2_TB2_CLKIO_N_6,
    input wire        mb1_FA2_TB2_CLKIO_N_2_mb1_FB2_TB2_CLKIO_N_4,
    input wire        mb1_FA2_TB2_CLKIO_N_3_mb1_FB2_TB2_CLKIO_N_3,
    input wire        mb1_FA2_TB2_CLKIO_N_4_mb1_FB2_TB2_CLKIO_N_2,
    input wire        mb1_FA2_TB2_CLKIO_N_5_mb1_FB2_TB2_IO_010,
    input wire        mb1_FA2_TB2_CLKIO_N_6_mb1_FB2_TB2_CLKIO_N_1,
    input wire        mb1_FA2_TB2_CLKIO_N_7_mb1_FB2_TB2_CLKIO_N_0,
    input wire        mb1_FA2_TB2_CLKIO_P_0_mb1_FB2_TB2_CLKIO_P_7,
    input wire        mb1_FA2_TB2_CLKIO_P_1_mb1_FB2_TB2_CLKIO_P_6,
    input wire        mb1_FA2_TB2_CLKIO_P_2_mb1_FB2_TB2_CLKIO_P_4,
    input wire        mb1_FA2_TB2_CLKIO_P_3_mb1_FB2_TB2_CLKIO_P_3,
    input wire        mb1_FA2_TB2_CLKIO_P_4_mb1_FB2_TB2_CLKIO_P_2,
    input wire        mb1_FA2_TB2_CLKIO_P_5_mb1_FB2_TB2_IO_011,
    input wire        mb1_FA2_TB2_CLKIO_P_6_mb1_FB2_TB2_CLKIO_P_1,
    input wire        mb1_FA2_TB2_CLKIO_P_7_mb1_FB2_TB2_CLKIO_P_0,
    input wire        mb1_FA2_TB2_IO_004_mb1_FB2_TB2_IO_006,
    input wire        mb1_FA2_TB2_IO_005_mb1_FB2_TB2_IO_007,
    input wire        mb1_FA2_TB2_IO_006_mb1_FB2_TB2_IO_004,
    input wire        mb1_FA2_TB2_IO_007_mb1_FB2_TB2_IO_005,
    input wire        mb1_FA2_TB2_IO_008_mb1_FB2_TB2_IO_022,
    input wire        mb1_FA2_TB2_IO_009_mb1_FB2_TB2_IO_023,
    input wire        mb1_FA2_TB2_IO_010_mb1_FB2_TB2_CLKIO_N_5,
    input wire        mb1_FA2_TB2_IO_011_mb1_FB2_TB2_CLKIO_P_5,
    input wire        mb1_FA2_TB2_IO_012_mb1_FB2_TB2_IO_012,
    input wire        mb1_FA2_TB2_IO_013_mb1_FB2_TB2_IO_013,
    input wire        mb1_FA2_TB2_IO_014_mb1_FB2_TB2_IO_016,
    input wire        mb1_FA2_TB2_IO_015_mb1_FB2_TB2_IO_017,
    input wire        mb1_FA2_TB2_IO_016_mb1_FB2_TB2_IO_014,
    input wire        mb1_FA2_TB2_IO_017_mb1_FB2_TB2_IO_015,
    input wire        mb1_FA2_TB2_IO_018_mb1_FB2_TB2_IO_032,
    input wire        mb1_FA2_TB2_IO_019_mb1_FB2_TB2_IO_033,
    input wire        mb1_FA2_TB2_IO_020_mb1_FB2_TB2_IO_030,
    input wire        mb1_FA2_TB2_IO_021_mb1_FB2_TB2_IO_031,
    input wire        mb1_FA2_TB2_IO_022_mb1_FB2_TB2_IO_008,
    input wire        mb1_FA2_TB2_IO_023_mb1_FB2_TB2_IO_009,
    input wire        mb1_FA2_TB2_IO_024_mb1_FB2_TB2_IO_026,
    input wire        mb1_FA2_TB2_IO_025_mb1_FB2_TB2_IO_027,
    input wire        mb1_FA2_TB2_IO_026_mb1_FB2_TB2_IO_024,
    input wire        mb1_FA2_TB2_IO_027_mb1_FB2_TB2_IO_025,
    input wire        mb1_FA2_TB2_IO_028_mb1_FB2_TB2_IO_042,
    input wire        mb1_FA2_TB2_IO_029_mb1_FB2_TB2_IO_043,
    input wire        mb1_FA2_TB2_IO_030_mb1_FB2_TB2_IO_020,
    input wire        mb1_FA2_TB2_IO_031_mb1_FB2_TB2_IO_021,
    input wire        mb1_FA2_TB2_IO_032_mb1_FB2_TB2_IO_018,
    input wire        mb1_FA2_TB2_IO_033_mb1_FB2_TB2_IO_019,
    input wire        mb1_FA2_TB2_IO_034_mb1_FB2_TB2_IO_036,
    input wire        mb1_FA2_TB2_IO_035_mb1_FB2_TB2_IO_037,
    input wire        mb1_FA2_TB2_IO_036_mb1_FB2_TB2_IO_034,
    input wire        mb1_FA2_TB2_IO_037_mb1_FB2_TB2_IO_035,
    input wire        mb1_FA2_TB2_IO_038_mb1_FB2_TB2_IO_052,
    input wire        mb1_FA2_TB2_IO_039_mb1_FB2_TB2_IO_053,
    input wire        mb1_FA2_TB2_IO_040_mb1_FB2_TB2_IO_050,
    input wire        mb1_FA2_TB2_IO_041_mb1_FB2_TB2_IO_051,
    input wire        mb1_FA2_TB2_IO_042_mb1_FB2_TB2_IO_028,
    input wire        mb1_FA2_TB2_IO_043_mb1_FB2_TB2_IO_029,
    input wire        mb1_FA2_TB2_IO_044_mb1_FB2_TB2_IO_046,
    input wire        mb1_FA2_TB2_IO_045_mb1_FB2_TB2_IO_047,
    input wire        mb1_FA2_TB2_IO_046_mb1_FB2_TB2_IO_044,
    input wire        mb1_FA2_TB2_IO_047_mb1_FB2_TB2_IO_045,
    input wire        mb1_FA2_TB2_IO_048_mb1_FB2_TB2_IO_062,
    input wire        mb1_FA2_TB2_IO_049_mb1_FB2_TB2_IO_063,
    input wire        mb1_FA2_TB2_IO_050_mb1_FB2_TB2_IO_040,
    input wire        mb1_FA2_TB2_IO_051_mb1_FB2_TB2_IO_041,
    input wire        mb1_FA2_TB2_IO_052_mb1_FB2_TB2_IO_038,
    input wire        mb1_FA2_TB2_IO_053_mb1_FB2_TB2_IO_039,
    input wire        mb1_FA2_TB2_IO_054_mb1_FB2_TB2_IO_056,
    input wire        mb1_FA2_TB2_IO_055_mb1_FB2_TB2_IO_057,
    input wire        mb1_FA2_TB2_IO_056_mb1_FB2_TB2_IO_054,
    input wire        mb1_FA2_TB2_IO_057_mb1_FB2_TB2_IO_055,
    input wire        mb1_FA2_TB2_IO_058_mb1_FB2_TB2_IO_072,
    input wire        mb1_FA2_TB2_IO_059_mb1_FB2_TB2_IO_073,
    input wire        mb1_FA2_TB2_IO_060_mb1_FB2_TB2_IO_070,
    input wire        mb1_FA2_TB2_IO_061_mb1_FB2_TB2_IO_071,
    input wire        mb1_FA2_TB2_IO_062_mb1_FB2_TB2_IO_048,
    input wire        mb1_FA2_TB2_IO_063_mb1_FB2_TB2_IO_049,
    input wire        mb1_FA2_TB2_IO_064_mb1_FB2_TB2_IO_066,
    input wire        mb1_FA2_TB2_IO_065_mb1_FB2_TB2_IO_067,
    input wire        mb1_FA2_TB2_IO_066_mb1_FB2_TB2_IO_064,
    input wire        mb1_FA2_TB2_IO_067_mb1_FB2_TB2_IO_065,
    input wire        mb1_FA2_TB2_IO_068_mb1_FB2_TB2_IO_082,
    input wire        mb1_FA2_TB2_IO_069_mb1_FB2_TB2_IO_083,
    input wire        mb1_FA2_TB2_IO_070_mb1_FB2_TB2_IO_060,
    input wire        mb1_FA2_TB2_IO_071_mb1_FB2_TB2_IO_061,
    input wire        mb1_FA2_TB2_IO_072_mb1_FB2_TB2_IO_058,
    input wire        mb1_FA2_TB2_IO_073_mb1_FB2_TB2_IO_059,
    input wire        mb1_FA2_TB2_IO_074_mb1_FB2_TB2_IO_076,
    input wire        mb1_FA2_TB2_IO_075_mb1_FB2_TB2_IO_077,
    input wire        mb1_FA2_TB2_IO_076_mb1_FB2_TB2_IO_074,
    input wire        mb1_FA2_TB2_IO_077_mb1_FB2_TB2_IO_075,
    input wire        mb1_FA2_TB2_IO_078_mb1_FB2_TB2_IO_092,
    input wire        mb1_FA2_TB2_IO_079_mb1_FB2_TB2_IO_093,
    input wire        mb1_FA2_TB2_IO_080_mb1_FB2_TB2_IO_090,
    input wire        mb1_FA2_TB2_IO_081_mb1_FB2_TB2_IO_091,
    input wire        mb1_FA2_TB2_IO_082_mb1_FB2_TB2_IO_068,
    input wire        mb1_FA2_TB2_IO_083_mb1_FB2_TB2_IO_069,
    input wire        mb1_FA2_TB2_IO_084_mb1_FB2_TB2_IO_086,
    input wire        mb1_FA2_TB2_IO_085_mb1_FB2_TB2_IO_087,
    input wire        mb1_FA2_TB2_IO_086_mb1_FB2_TB2_IO_084,
    input wire        mb1_FA2_TB2_IO_087_mb1_FB2_TB2_IO_085,
    input wire        mb1_FA2_TB2_IO_088_mb1_FB2_TB2_IO_102,
    input wire        mb1_FA2_TB2_IO_089_mb1_FB2_TB2_IO_103,
    input wire        mb1_FA2_TB2_IO_090_mb1_FB2_TB2_IO_080,
    input wire        mb1_FA2_TB2_IO_091_mb1_FB2_TB2_IO_081,
    input wire        mb1_FA2_TB2_IO_092_mb1_FB2_TB2_IO_078,
    input wire        mb1_FA2_TB2_IO_093_mb1_FB2_TB2_IO_079,
    input wire        mb1_FA2_TB2_IO_094_mb1_FB2_TB2_IO_096,
    input wire        mb1_FA2_TB2_IO_095_mb1_FB2_TB2_IO_097,
    input wire        mb1_FA2_TB2_IO_096_mb1_FB2_TB2_IO_094,
    input wire        mb1_FA2_TB2_IO_097_mb1_FB2_TB2_IO_095,
    input wire        mb1_FA2_TB2_IO_098_mb1_FB2_TB2_IO_112,
    input wire        mb1_FA2_TB2_IO_099_mb1_FB2_TB2_IO_113,
    input wire        mb1_FA2_TB2_IO_100_mb1_FB2_TB2_IO_110,
    input wire        mb1_FA2_TB2_IO_101_mb1_FB2_TB2_IO_111,
    input wire        mb1_FA2_TB2_IO_102_mb1_FB2_TB2_IO_088,
    input wire        mb1_FA2_TB2_IO_103_mb1_FB2_TB2_IO_089,
    input wire        mb1_FA2_TB2_IO_104_mb1_FB2_TB2_IO_106,
    input wire        mb1_FA2_TB2_IO_105_mb1_FB2_TB2_IO_107,
    input wire        mb1_FA2_TB2_IO_106_mb1_FB2_TB2_IO_104,
    input wire        mb1_FA2_TB2_IO_107_mb1_FB2_TB2_IO_105,
    input wire        mb1_FA2_TB2_IO_108_mb1_FB2_TB2_IO_122,
    input wire        mb1_FA2_TB2_IO_109_mb1_FB2_TB2_IO_123,
    input wire        mb1_FA2_TB2_IO_110_mb1_FB2_TB2_IO_100,
    input wire        mb1_FA2_TB2_IO_111_mb1_FB2_TB2_IO_101,
    input wire        mb1_FA2_TB2_IO_112_mb1_FB2_TB2_IO_098,
    input wire        mb1_FA2_TB2_IO_113_mb1_FB2_TB2_IO_099,
    input wire        mb1_FA2_TB2_IO_114_mb1_FB2_TB2_IO_116,
    input wire        mb1_FA2_TB2_IO_115_mb1_FB2_TB2_IO_117,
    input wire        mb1_FA2_TB2_IO_116_mb1_FB2_TB2_IO_114,
    input wire        mb1_FA2_TB2_IO_117_mb1_FB2_TB2_IO_115,
    input wire        mb1_FA2_TB2_IO_118_mb1_FB2_TB2_IO_132,
    input wire        mb1_FA2_TB2_IO_119_mb1_FB2_TB2_IO_133,
    input wire        mb1_FA2_TB2_IO_120_mb1_FB2_TB2_IO_130,
    input wire        mb1_FA2_TB2_IO_121_mb1_FB2_TB2_IO_131,
    input wire        mb1_FA2_TB2_IO_122_mb1_FB2_TB2_IO_108,
    input wire        mb1_FA2_TB2_IO_123_mb1_FB2_TB2_IO_109,
    input wire        mb1_FA2_TB2_IO_124_mb1_FB2_TB2_IO_126,
    input wire        mb1_FA2_TB2_IO_125_mb1_FB2_TB2_IO_127,
    input wire        mb1_FA2_TB2_IO_126_mb1_FB2_TB2_IO_124,
    input wire        mb1_FA2_TB2_IO_127_mb1_FB2_TB2_IO_125,
    input wire        mb1_FA2_TB2_IO_130_mb1_FB2_TB2_IO_120,
    input wire        mb1_FA2_TB2_IO_131_mb1_FB2_TB2_IO_121,
    input wire        mb1_FA2_TB2_IO_132_mb1_FB2_TB2_IO_118,
    input wire        mb1_FA2_TB2_IO_133_mb1_FB2_TB2_IO_119,
    input wire        mb1_FA2_TB2_IO_134_mb1_FB2_TB2_IO_136,
    input wire        mb1_FA2_TB2_IO_136_mb1_FB2_TB2_IO_134,
    input wire        mb1_FA2_TA1_CLKIO_N_0_mb1_FB2_BA0_CLKIO_N_7,
    input wire        mb1_FA2_TA1_CLKIO_N_1_mb1_FB2_BA0_CLKIO_N_6,
    input wire        mb1_FA2_TA1_CLKIO_N_2_mb1_FB2_BA0_CLKIO_N_4,
    input wire        mb1_FA2_TA1_CLKIO_N_3_mb1_FB2_BA0_CLKIO_N_3,
    input wire        mb1_FA2_TA1_CLKIO_N_4_mb1_FB2_BA0_CLKIO_N_2,
    input wire        mb1_FA2_TA1_CLKIO_N_5_mb1_FB2_BA0_IO_010,
    input wire        mb1_FA2_TA1_CLKIO_N_6_mb1_FB2_BA0_CLKIO_N_1,
    input wire        mb1_FA2_TA1_CLKIO_N_7_mb1_FB2_BA0_CLKIO_N_0,
    input wire        mb1_FA2_TA1_CLKIO_P_0_mb1_FB2_BA0_CLKIO_P_7,
    input wire        mb1_FA2_TA1_CLKIO_P_1_mb1_FB2_BA0_CLKIO_P_6,
    input wire        mb1_FA2_TA1_CLKIO_P_2_mb1_FB2_BA0_CLKIO_P_4,
    input wire        mb1_FA2_TA1_CLKIO_P_3_mb1_FB2_BA0_CLKIO_P_3,
    input wire        mb1_FA2_TA1_CLKIO_P_4_mb1_FB2_BA0_CLKIO_P_2,
    input wire        mb1_FA2_TA1_CLKIO_P_5_mb1_FB2_BA0_IO_011,
    input wire        mb1_FA2_TA1_CLKIO_P_6_mb1_FB2_BA0_CLKIO_P_1,
    input wire        mb1_FA2_TA1_CLKIO_P_7_mb1_FB2_BA0_CLKIO_P_0,
    input wire        mb1_FA2_TA1_IO_004_mb1_FB2_BA0_IO_006,
    input wire        mb1_FA2_TA1_IO_005_mb1_FB2_BA0_IO_007,
    input wire        mb1_FA2_TA1_IO_006_mb1_FB2_BA0_IO_004,
    input wire        mb1_FA2_TA1_IO_007_mb1_FB2_BA0_IO_005,
    input wire        mb1_FA2_TA1_IO_008_mb1_FB2_BA0_IO_022,
    input wire        mb1_FA2_TA1_IO_009_mb1_FB2_BA0_IO_023,
    input wire        mb1_FA2_TA1_IO_010_mb1_FB2_BA0_CLKIO_N_5,
    input wire        mb1_FA2_TA1_IO_011_mb1_FB2_BA0_CLKIO_P_5,
    input wire        mb1_FA2_TA1_IO_012_mb1_FB2_BA0_IO_012,
    input wire        mb1_FA2_TA1_IO_013_mb1_FB2_BA0_IO_013,
    input wire        mb1_FA2_TA1_IO_014_mb1_FB2_BA0_IO_016,
    input wire        mb1_FA2_TA1_IO_015_mb1_FB2_BA0_IO_017,
    input wire        mb1_FA2_TA1_IO_016_mb1_FB2_BA0_IO_014,
    input wire        mb1_FA2_TA1_IO_017_mb1_FB2_BA0_IO_015,
    input wire        mb1_FA2_TA1_IO_018_mb1_FB2_BA0_IO_032,
    input wire        mb1_FA2_TA1_IO_019_mb1_FB2_BA0_IO_033,
    input wire        mb1_FA2_TA1_IO_020_mb1_FB2_BA0_IO_030,
    input wire        mb1_FA2_TA1_IO_021_mb1_FB2_BA0_IO_031,
    input wire        mb1_FA2_TA1_IO_022_mb1_FB2_BA0_IO_008,
    input wire        mb1_FA2_TA1_IO_023_mb1_FB2_BA0_IO_009,
    input wire        mb1_FA2_TA1_IO_024_mb1_FB2_BA0_IO_026,
    input wire        mb1_FA2_TA1_IO_025_mb1_FB2_BA0_IO_027,
    input wire        mb1_FA2_TA1_IO_026_mb1_FB2_BA0_IO_024,
    input wire        mb1_FA2_TA1_IO_027_mb1_FB2_BA0_IO_025,
    input wire        mb1_FA2_TA1_IO_028_mb1_FB2_BA0_IO_042,
    input wire        mb1_FA2_TA1_IO_029_mb1_FB2_BA0_IO_043,
    input wire        mb1_FA2_TA1_IO_030_mb1_FB2_BA0_IO_020,
    input wire        mb1_FA2_TA1_IO_031_mb1_FB2_BA0_IO_021,
    input wire        mb1_FA2_TA1_IO_032_mb1_FB2_BA0_IO_018,
    input wire        mb1_FA2_TA1_IO_033_mb1_FB2_BA0_IO_019,
    input wire        mb1_FA2_TA1_IO_034_mb1_FB2_BA0_IO_036,
    input wire        mb1_FA2_TA1_IO_035_mb1_FB2_BA0_IO_037,
    input wire        mb1_FA2_TA1_IO_036_mb1_FB2_BA0_IO_034,
    input wire        mb1_FA2_TA1_IO_037_mb1_FB2_BA0_IO_035,
    input wire        mb1_FA2_TA1_IO_038_mb1_FB2_BA0_IO_052,
    input wire        mb1_FA2_TA1_IO_039_mb1_FB2_BA0_IO_053,
    input wire        mb1_FA2_TA1_IO_040_mb1_FB2_BA0_IO_050,
    input wire        mb1_FA2_TA1_IO_041_mb1_FB2_BA0_IO_051,
    input wire        mb1_FA2_TA1_IO_042_mb1_FB2_BA0_IO_028,
    input wire        mb1_FA2_TA1_IO_043_mb1_FB2_BA0_IO_029,
    input wire        mb1_FA2_TA1_IO_044_mb1_FB2_BA0_IO_046,
    input wire        mb1_FA2_TA1_IO_045_mb1_FB2_BA0_IO_047,
    input wire        mb1_FA2_TA1_IO_046_mb1_FB2_BA0_IO_044,
    input wire        mb1_FA2_TA1_IO_047_mb1_FB2_BA0_IO_045,
    input wire        mb1_FA2_TA1_IO_048_mb1_FB2_BA0_IO_062,
    input wire        mb1_FA2_TA1_IO_049_mb1_FB2_BA0_IO_063,
    input wire        mb1_FA2_TA1_IO_050_mb1_FB2_BA0_IO_040,
    input wire        mb1_FA2_TA1_IO_051_mb1_FB2_BA0_IO_041,
    input wire        mb1_FA2_TA1_IO_052_mb1_FB2_BA0_IO_038,
    input wire        mb1_FA2_TA1_IO_053_mb1_FB2_BA0_IO_039,
    input wire        mb1_FA2_TA1_IO_054_mb1_FB2_BA0_IO_056,
    input wire        mb1_FA2_TA1_IO_055_mb1_FB2_BA0_IO_057,
    input wire        mb1_FA2_TA1_IO_056_mb1_FB2_BA0_IO_054,
    input wire        mb1_FA2_TA1_IO_057_mb1_FB2_BA0_IO_055,
    input wire        mb1_FA2_TA1_IO_058_mb1_FB2_BA0_IO_072,
    input wire        mb1_FA2_TA1_IO_059_mb1_FB2_BA0_IO_073,
    input wire        mb1_FA2_TA1_IO_060_mb1_FB2_BA0_IO_070,
    input wire        mb1_FA2_TA1_IO_061_mb1_FB2_BA0_IO_071,
    input wire        mb1_FA2_TA1_IO_062_mb1_FB2_BA0_IO_048,
    input wire        mb1_FA2_TA1_IO_063_mb1_FB2_BA0_IO_049,
    input wire        mb1_FA2_TA1_IO_064_mb1_FB2_BA0_IO_066,
    input wire        mb1_FA2_TA1_IO_065_mb1_FB2_BA0_IO_067,
    input wire        mb1_FA2_TA1_IO_066_mb1_FB2_BA0_IO_064,
    input wire        mb1_FA2_TA1_IO_067_mb1_FB2_BA0_IO_065,
    input wire        mb1_FA2_TA1_IO_068_mb1_FB2_BA0_IO_082,
    input wire        mb1_FA2_TA1_IO_069_mb1_FB2_BA0_IO_083,
    input wire        mb1_FA2_TA1_IO_070_mb1_FB2_BA0_IO_060,
    input wire        mb1_FA2_TA1_IO_071_mb1_FB2_BA0_IO_061,
    input wire        mb1_FA2_TA1_IO_072_mb1_FB2_BA0_IO_058,
    input wire        mb1_FA2_TA1_IO_073_mb1_FB2_BA0_IO_059,
    input wire        mb1_FA2_TA1_IO_074_mb1_FB2_BA0_IO_076,
    input wire        mb1_FA2_TA1_IO_075_mb1_FB2_BA0_IO_077,
    input wire        mb1_FA2_TA1_IO_076_mb1_FB2_BA0_IO_074,
    input wire        mb1_FA2_TA1_IO_077_mb1_FB2_BA0_IO_075,
    input wire        mb1_FA2_TA1_IO_078_mb1_FB2_BA0_IO_092,
    input wire        mb1_FA2_TA1_IO_079_mb1_FB2_BA0_IO_093,
    input wire        mb1_FA2_TA1_IO_080_mb1_FB2_BA0_IO_090,
    input wire        mb1_FA2_TA1_IO_081_mb1_FB2_BA0_IO_091,
    input wire        mb1_FA2_TA1_IO_082_mb1_FB2_BA0_IO_068,
    input wire        mb1_FA2_TA1_IO_083_mb1_FB2_BA0_IO_069,
    input wire        mb1_FA2_TA1_IO_084_mb1_FB2_BA0_IO_086,
    input wire        mb1_FA2_TA1_IO_085_mb1_FB2_BA0_IO_087,
    input wire        mb1_FA2_TA1_IO_086_mb1_FB2_BA0_IO_084,
    input wire        mb1_FA2_TA1_IO_087_mb1_FB2_BA0_IO_085,
    input wire        mb1_FA2_TA1_IO_088_mb1_FB2_BA0_IO_102,
    input wire        mb1_FA2_TA1_IO_089_mb1_FB2_BA0_IO_103,
    input wire        mb1_FA2_TA1_IO_090_mb1_FB2_BA0_IO_080,
    input wire        mb1_FA2_TA1_IO_091_mb1_FB2_BA0_IO_081,
    input wire        mb1_FA2_TA1_IO_092_mb1_FB2_BA0_IO_078,
    input wire        mb1_FA2_TA1_IO_093_mb1_FB2_BA0_IO_079,
    input wire        mb1_FA2_TA1_IO_094_mb1_FB2_BA0_IO_096,
    input wire        mb1_FA2_TA1_IO_095_mb1_FB2_BA0_IO_097,
    input wire        mb1_FA2_TA1_IO_096_mb1_FB2_BA0_IO_094,
    input wire        mb1_FA2_TA1_IO_097_mb1_FB2_BA0_IO_095,
    input wire        mb1_FA2_TA1_IO_098_mb1_FB2_BA0_IO_112,
    input wire        mb1_FA2_TA1_IO_099_mb1_FB2_BA0_IO_113,
    input wire        mb1_FA2_TA1_IO_100_mb1_FB2_BA0_IO_110,
    input wire        mb1_FA2_TA1_IO_101_mb1_FB2_BA0_IO_111,
    input wire        mb1_FA2_TA1_IO_102_mb1_FB2_BA0_IO_088,
    input wire        mb1_FA2_TA1_IO_103_mb1_FB2_BA0_IO_089,
    input wire        mb1_FA2_TA1_IO_104_mb1_FB2_BA0_IO_106,
    input wire        mb1_FA2_TA1_IO_105_mb1_FB2_BA0_IO_107,
    input wire        mb1_FA2_TA1_IO_106_mb1_FB2_BA0_IO_104,
    input wire        mb1_FA2_TA1_IO_107_mb1_FB2_BA0_IO_105,
    input wire        mb1_FA2_TA1_IO_108_mb1_FB2_BA0_IO_122,
    input wire        mb1_FA2_TA1_IO_109_mb1_FB2_BA0_IO_123,
    input wire        mb1_FA2_TA1_IO_110_mb1_FB2_BA0_IO_100,
    input wire        mb1_FA2_TA1_IO_111_mb1_FB2_BA0_IO_101,
    input wire        mb1_FA2_TA1_IO_112_mb1_FB2_BA0_IO_098,
    input wire        mb1_FA2_TA1_IO_113_mb1_FB2_BA0_IO_099,
    input wire        mb1_FA2_TA1_IO_114_mb1_FB2_BA0_IO_116,
    input wire        mb1_FA2_TA1_IO_115_mb1_FB2_BA0_IO_117,
    input wire        mb1_FA2_TA1_IO_116_mb1_FB2_BA0_IO_114,
    input wire        mb1_FA2_TA1_IO_117_mb1_FB2_BA0_IO_115,
    input wire        mb1_FA2_TA1_IO_118_mb1_FB2_BA0_IO_132,
    input wire        mb1_FA2_TA1_IO_119_mb1_FB2_BA0_IO_133,
    input wire        mb1_FA2_TA1_IO_120_mb1_FB2_BA0_IO_130,
    input wire        mb1_FA2_TA1_IO_121_mb1_FB2_BA0_IO_131,
    input wire        mb1_FA2_TA1_IO_122_mb1_FB2_BA0_IO_108,
    input wire        mb1_FA2_TA1_IO_123_mb1_FB2_BA0_IO_109,
    input wire        mb1_FA2_TA1_IO_124_mb1_FB2_BA0_IO_126,
    input wire        mb1_FA2_TA1_IO_125_mb1_FB2_BA0_IO_127,
    input wire        mb1_FA2_TA1_IO_126_mb1_FB2_BA0_IO_124,
    input wire        mb1_FA2_TA1_IO_127_mb1_FB2_BA0_IO_125,
    input wire        mb1_FA2_TA1_IO_130_mb1_FB2_BA0_IO_120,
    input wire        mb1_FA2_TA1_IO_131_mb1_FB2_BA0_IO_121,
    input wire        mb1_FA2_TA1_IO_132_mb1_FB2_BA0_IO_118,
    input wire        mb1_FA2_TA1_IO_133_mb1_FB2_BA0_IO_119,
    input wire        mb1_FA2_TA1_IO_134_mb1_FB2_BA0_IO_136,
    input wire        mb1_FA2_TA1_IO_136_mb1_FB2_BA0_IO_134,
    input wire        mb1_FA2_BB0_CLKIO_N_0_mb1_FB2_BA1_CLKIO_N_7,
    input wire        mb1_FA2_BB0_CLKIO_N_1_mb1_FB2_BA1_CLKIO_N_6,
    input wire        mb1_FA2_BB0_CLKIO_N_2_mb1_FB2_BA1_CLKIO_N_4,
    input wire        mb1_FA2_BB0_CLKIO_N_3_mb1_FB2_BA1_CLKIO_N_3,
    input wire        mb1_FA2_BB0_CLKIO_N_4_mb1_FB2_BA1_CLKIO_N_2,
    input wire        mb1_FA2_BB0_CLKIO_N_5_mb1_FB2_BA1_IO_010,
    input wire        mb1_FA2_BB0_CLKIO_N_6_mb1_FB2_BA1_CLKIO_N_1,
    input wire        mb1_FA2_BB0_CLKIO_N_7_mb1_FB2_BA1_CLKIO_N_0,
    input wire        mb1_FA2_BB0_CLKIO_P_0_mb1_FB2_BA1_CLKIO_P_7,
    input wire        mb1_FA2_BB0_CLKIO_P_1_mb1_FB2_BA1_CLKIO_P_6,
    input wire        mb1_FA2_BB0_CLKIO_P_2_mb1_FB2_BA1_CLKIO_P_4,
    input wire        mb1_FA2_BB0_CLKIO_P_3_mb1_FB2_BA1_CLKIO_P_3,
    input wire        mb1_FA2_BB0_CLKIO_P_4_mb1_FB2_BA1_CLKIO_P_2,
    input wire        mb1_FA2_BB0_CLKIO_P_5_mb1_FB2_BA1_IO_011,
    input wire        mb1_FA2_BB0_CLKIO_P_6_mb1_FB2_BA1_CLKIO_P_1,
    input wire        mb1_FA2_BB0_CLKIO_P_7_mb1_FB2_BA1_CLKIO_P_0,
    input wire        mb1_FA2_BB0_IO_004_mb1_FB2_BA1_IO_006,
    input wire        mb1_FA2_BB0_IO_005_mb1_FB2_BA1_IO_007,
    input wire        mb1_FA2_BB0_IO_006_mb1_FB2_BA1_IO_004,
    input wire        mb1_FA2_BB0_IO_007_mb1_FB2_BA1_IO_005,
    input wire        mb1_FA2_BB0_IO_008_mb1_FB2_BA1_IO_022,
    input wire        mb1_FA2_BB0_IO_009_mb1_FB2_BA1_IO_023,
    input wire        mb1_FA2_BB0_IO_010_mb1_FB2_BA1_CLKIO_N_5,
    input wire        mb1_FA2_BB0_IO_011_mb1_FB2_BA1_CLKIO_P_5,
    input wire        mb1_FA2_BB0_IO_012_mb1_FB2_BA1_IO_012,
    input wire        mb1_FA2_BB0_IO_013_mb1_FB2_BA1_IO_013,
    input wire        mb1_FA2_BB0_IO_014_mb1_FB2_BA1_IO_016,
    input wire        mb1_FA2_BB0_IO_015_mb1_FB2_BA1_IO_017,
    input wire        mb1_FA2_BB0_IO_016_mb1_FB2_BA1_IO_014,
    input wire        mb1_FA2_BB0_IO_017_mb1_FB2_BA1_IO_015,
    input wire        mb1_FA2_BB0_IO_018_mb1_FB2_BA1_IO_032,
    input wire        mb1_FA2_BB0_IO_019_mb1_FB2_BA1_IO_033,
    input wire        mb1_FA2_BB0_IO_020_mb1_FB2_BA1_IO_030,
    input wire        mb1_FA2_BB0_IO_021_mb1_FB2_BA1_IO_031,
    input wire        mb1_FA2_BB0_IO_022_mb1_FB2_BA1_IO_008,
    input wire        mb1_FA2_BB0_IO_023_mb1_FB2_BA1_IO_009,
    input wire        mb1_FA2_BB0_IO_024_mb1_FB2_BA1_IO_026,
    input wire        mb1_FA2_BB0_IO_025_mb1_FB2_BA1_IO_027,
    input wire        mb1_FA2_BB0_IO_026_mb1_FB2_BA1_IO_024,
    input wire        mb1_FA2_BB0_IO_027_mb1_FB2_BA1_IO_025,
    input wire        mb1_FA2_BB0_IO_028_mb1_FB2_BA1_IO_042,
    input wire        mb1_FA2_BB0_IO_029_mb1_FB2_BA1_IO_043,
    input wire        mb1_FA2_BB0_IO_030_mb1_FB2_BA1_IO_020,
    input wire        mb1_FA2_BB0_IO_031_mb1_FB2_BA1_IO_021,
    input wire        mb1_FA2_BB0_IO_032_mb1_FB2_BA1_IO_018,
    input wire        mb1_FA2_BB0_IO_033_mb1_FB2_BA1_IO_019,
    input wire        mb1_FA2_BB0_IO_034_mb1_FB2_BA1_IO_036,
    input wire        mb1_FA2_BB0_IO_035_mb1_FB2_BA1_IO_037,
    input wire        mb1_FA2_BB0_IO_036_mb1_FB2_BA1_IO_034,
    input wire        mb1_FA2_BB0_IO_037_mb1_FB2_BA1_IO_035,
    input wire        mb1_FA2_BB0_IO_038_mb1_FB2_BA1_IO_052,
    input wire        mb1_FA2_BB0_IO_039_mb1_FB2_BA1_IO_053,
    input wire        mb1_FA2_BB0_IO_040_mb1_FB2_BA1_IO_050,
    input wire        mb1_FA2_BB0_IO_041_mb1_FB2_BA1_IO_051,
    input wire        mb1_FA2_BB0_IO_042_mb1_FB2_BA1_IO_028,
    input wire        mb1_FA2_BB0_IO_043_mb1_FB2_BA1_IO_029,
    input wire        mb1_FA2_BB0_IO_044_mb1_FB2_BA1_IO_046,
    input wire        mb1_FA2_BB0_IO_045_mb1_FB2_BA1_IO_047,
    input wire        mb1_FA2_BB0_IO_046_mb1_FB2_BA1_IO_044,
    input wire        mb1_FA2_BB0_IO_047_mb1_FB2_BA1_IO_045,
    input wire        mb1_FA2_BB0_IO_048_mb1_FB2_BA1_IO_062,
    input wire        mb1_FA2_BB0_IO_049_mb1_FB2_BA1_IO_063,
    input wire        mb1_FA2_BB0_IO_050_mb1_FB2_BA1_IO_040,
    input wire        mb1_FA2_BB0_IO_051_mb1_FB2_BA1_IO_041,
    input wire        mb1_FA2_BB0_IO_052_mb1_FB2_BA1_IO_038,
    input wire        mb1_FA2_BB0_IO_053_mb1_FB2_BA1_IO_039,
    input wire        mb1_FA2_BB0_IO_054_mb1_FB2_BA1_IO_056,
    input wire        mb1_FA2_BB0_IO_055_mb1_FB2_BA1_IO_057,
    input wire        mb1_FA2_BB0_IO_056_mb1_FB2_BA1_IO_054,
    input wire        mb1_FA2_BB0_IO_057_mb1_FB2_BA1_IO_055,
    input wire        mb1_FA2_BB0_IO_058_mb1_FB2_BA1_IO_072,
    input wire        mb1_FA2_BB0_IO_059_mb1_FB2_BA1_IO_073,
    input wire        mb1_FA2_BB0_IO_060_mb1_FB2_BA1_IO_070,
    input wire        mb1_FA2_BB0_IO_061_mb1_FB2_BA1_IO_071,
    input wire        mb1_FA2_BB0_IO_062_mb1_FB2_BA1_IO_048,
    input wire        mb1_FA2_BB0_IO_063_mb1_FB2_BA1_IO_049,
    input wire        mb1_FA2_BB0_IO_064_mb1_FB2_BA1_IO_066,
    input wire        mb1_FA2_BB0_IO_065_mb1_FB2_BA1_IO_067,
    input wire        mb1_FA2_BB0_IO_066_mb1_FB2_BA1_IO_064,
    input wire        mb1_FA2_BB0_IO_067_mb1_FB2_BA1_IO_065,
    input wire        mb1_FA2_BB0_IO_068_mb1_FB2_BA1_IO_082,
    input wire        mb1_FA2_BB0_IO_069_mb1_FB2_BA1_IO_083,
    input wire        mb1_FA2_BB0_IO_070_mb1_FB2_BA1_IO_060,
    input wire        mb1_FA2_BB0_IO_071_mb1_FB2_BA1_IO_061,
    input wire        mb1_FA2_BB0_IO_072_mb1_FB2_BA1_IO_058,
    input wire        mb1_FA2_BB0_IO_073_mb1_FB2_BA1_IO_059,
    input wire        mb1_FA2_BB0_IO_074_mb1_FB2_BA1_IO_076,
    input wire        mb1_FA2_BB0_IO_075_mb1_FB2_BA1_IO_077,
    input wire        mb1_FA2_BB0_IO_076_mb1_FB2_BA1_IO_074,
    input wire        mb1_FA2_BB0_IO_077_mb1_FB2_BA1_IO_075,
    input wire        mb1_FA2_BB0_IO_078_mb1_FB2_BA1_IO_092,
    input wire        mb1_FA2_BB0_IO_079_mb1_FB2_BA1_IO_093,
    input wire        mb1_FA2_BB0_IO_080_mb1_FB2_BA1_IO_090,
    input wire        mb1_FA2_BB0_IO_081_mb1_FB2_BA1_IO_091,
    input wire        mb1_FA2_BB0_IO_082_mb1_FB2_BA1_IO_068,
    input wire        mb1_FA2_BB0_IO_083_mb1_FB2_BA1_IO_069,
    input wire        mb1_FA2_BB0_IO_084_mb1_FB2_BA1_IO_086,
    input wire        mb1_FA2_BB0_IO_085_mb1_FB2_BA1_IO_087,
    input wire        mb1_FA2_BB0_IO_086_mb1_FB2_BA1_IO_084,
    input wire        mb1_FA2_BB0_IO_087_mb1_FB2_BA1_IO_085,
    input wire        mb1_FA2_BB0_IO_088_mb1_FB2_BA1_IO_102,
    input wire        mb1_FA2_BB0_IO_089_mb1_FB2_BA1_IO_103,
    input wire        mb1_FA2_BB0_IO_090_mb1_FB2_BA1_IO_080,
    input wire        mb1_FA2_BB0_IO_091_mb1_FB2_BA1_IO_081,
    input wire        mb1_FA2_BB0_IO_092_mb1_FB2_BA1_IO_078,
    input wire        mb1_FA2_BB0_IO_093_mb1_FB2_BA1_IO_079,
    input wire        mb1_FA2_BB0_IO_094_mb1_FB2_BA1_IO_096,
    input wire        mb1_FA2_BB0_IO_095_mb1_FB2_BA1_IO_097,
    input wire        mb1_FA2_BB0_IO_096_mb1_FB2_BA1_IO_094,
    input wire        mb1_FA2_BB0_IO_097_mb1_FB2_BA1_IO_095,
    input wire        mb1_FA2_BB0_IO_098_mb1_FB2_BA1_IO_112,
    input wire        mb1_FA2_BB0_IO_099_mb1_FB2_BA1_IO_113,
    input wire        mb1_FA2_BB0_IO_100_mb1_FB2_BA1_IO_110,
    input wire        mb1_FA2_BB0_IO_101_mb1_FB2_BA1_IO_111,
    input wire        mb1_FA2_BB0_IO_102_mb1_FB2_BA1_IO_088,
    input wire        mb1_FA2_BB0_IO_103_mb1_FB2_BA1_IO_089,
    input wire        mb1_FA2_BB0_IO_104_mb1_FB2_BA1_IO_106,
    input wire        mb1_FA2_BB0_IO_105_mb1_FB2_BA1_IO_107,
    input wire        mb1_FA2_BB0_IO_106_mb1_FB2_BA1_IO_104,
    input wire        mb1_FA2_BB0_IO_107_mb1_FB2_BA1_IO_105,
    input wire        mb1_FA2_BB0_IO_108_mb1_FB2_BA1_IO_122,
    input wire        mb1_FA2_BB0_IO_109_mb1_FB2_BA1_IO_123,
    input wire        mb1_FA2_BB0_IO_110_mb1_FB2_BA1_IO_100,
    input wire        mb1_FA2_BB0_IO_111_mb1_FB2_BA1_IO_101,
    input wire        mb1_FA2_BB0_IO_112_mb1_FB2_BA1_IO_098,
    input wire        mb1_FA2_BB0_IO_113_mb1_FB2_BA1_IO_099,
    input wire        mb1_FA2_BB0_IO_114_mb1_FB2_BA1_IO_116,
    input wire        mb1_FA2_BB0_IO_115_mb1_FB2_BA1_IO_117,
    input wire        mb1_FA2_BB0_IO_116_mb1_FB2_BA1_IO_114,
    input wire        mb1_FA2_BB0_IO_117_mb1_FB2_BA1_IO_115,
    input wire        mb1_FA2_BB0_IO_118_mb1_FB2_BA1_IO_132,
    input wire        mb1_FA2_BB0_IO_119_mb1_FB2_BA1_IO_133,
    input wire        mb1_FA2_BB0_IO_120_mb1_FB2_BA1_IO_130,
    input wire        mb1_FA2_BB0_IO_121_mb1_FB2_BA1_IO_131,
    input wire        mb1_FA2_BB0_IO_122_mb1_FB2_BA1_IO_108,
    input wire        mb1_FA2_BB0_IO_123_mb1_FB2_BA1_IO_109,
    input wire        mb1_FA2_BB0_IO_124_mb1_FB2_BA1_IO_126,
    input wire        mb1_FA2_BB0_IO_125_mb1_FB2_BA1_IO_127,
    input wire        mb1_FA2_BB0_IO_126_mb1_FB2_BA1_IO_124,
    input wire        mb1_FA2_BB0_IO_127_mb1_FB2_BA1_IO_125,
    input wire        mb1_FA2_BB0_IO_130_mb1_FB2_BA1_IO_120,
    input wire        mb1_FA2_BB0_IO_131_mb1_FB2_BA1_IO_121,
    input wire        mb1_FA2_BB0_IO_132_mb1_FB2_BA1_IO_118,
    input wire        mb1_FA2_BB0_IO_133_mb1_FB2_BA1_IO_119,
    input wire        mb1_FA2_BB0_IO_134_mb1_FB2_BA1_IO_136,
    input wire        mb1_FA2_BB0_IO_136_mb1_FB2_BA1_IO_134,
    input wire        mb1_FA2_BA2_CLKIO_N_0_mb1_FB2_BA2_CLKIO_N_7,
    input wire        mb1_FA2_BA2_CLKIO_N_1_mb1_FB2_BA2_CLKIO_N_6,
    input wire        mb1_FA2_BA2_CLKIO_N_2_mb1_FB2_BA2_CLKIO_N_4,
    input wire        mb1_FA2_BA2_CLKIO_N_3_mb1_FB2_BA2_CLKIO_N_3,
    input wire        mb1_FA2_BA2_CLKIO_N_4_mb1_FB2_BA2_CLKIO_N_2,
    input wire        mb1_FA2_BA2_CLKIO_N_5_mb1_FB2_BA2_IO_010,
    input wire        mb1_FA2_BA2_CLKIO_N_6_mb1_FB2_BA2_CLKIO_N_1,
    input wire        mb1_FA2_BA2_CLKIO_N_7_mb1_FB2_BA2_CLKIO_N_0,
    input wire        mb1_FA2_BA2_CLKIO_P_0_mb1_FB2_BA2_CLKIO_P_7,
    input wire        mb1_FA2_BA2_CLKIO_P_1_mb1_FB2_BA2_CLKIO_P_6,
    input wire        mb1_FA2_BA2_CLKIO_P_2_mb1_FB2_BA2_CLKIO_P_4,
    input wire        mb1_FA2_BA2_CLKIO_P_3_mb1_FB2_BA2_CLKIO_P_3,
    input wire        mb1_FA2_BA2_CLKIO_P_4_mb1_FB2_BA2_CLKIO_P_2,
    input wire        mb1_FA2_BA2_CLKIO_P_5_mb1_FB2_BA2_IO_011,
    input wire        mb1_FA2_BA2_CLKIO_P_6_mb1_FB2_BA2_CLKIO_P_1,
    input wire        mb1_FA2_BA2_CLKIO_P_7_mb1_FB2_BA2_CLKIO_P_0,
    input wire        mb1_FA2_BA2_IO_004_mb1_FB2_BA2_IO_006,
    input wire        mb1_FA2_BA2_IO_005_mb1_FB2_BA2_IO_007,
    input wire        mb1_FA2_BA2_IO_006_mb1_FB2_BA2_IO_004,
    input wire        mb1_FA2_BA2_IO_007_mb1_FB2_BA2_IO_005,
    input wire        mb1_FA2_BA2_IO_008_mb1_FB2_BA2_IO_022,
    input wire        mb1_FA2_BA2_IO_009_mb1_FB2_BA2_IO_023,
    input wire        mb1_FA2_BA2_IO_010_mb1_FB2_BA2_CLKIO_N_5,
    input wire        mb1_FA2_BA2_IO_011_mb1_FB2_BA2_CLKIO_P_5,
    input wire        mb1_FA2_BA2_IO_012_mb1_FB2_BA2_IO_012,
    input wire        mb1_FA2_BA2_IO_013_mb1_FB2_BA2_IO_013,
    input wire        mb1_FA2_BA2_IO_014_mb1_FB2_BA2_IO_016,
    input wire        mb1_FA2_BA2_IO_015_mb1_FB2_BA2_IO_017,
    input wire        mb1_FA2_BA2_IO_016_mb1_FB2_BA2_IO_014,
    input wire        mb1_FA2_BA2_IO_017_mb1_FB2_BA2_IO_015,
    input wire        mb1_FA2_BA2_IO_018_mb1_FB2_BA2_IO_032,
    input wire        mb1_FA2_BA2_IO_019_mb1_FB2_BA2_IO_033,
    input wire        mb1_FA2_BA2_IO_020_mb1_FB2_BA2_IO_030,
    input wire        mb1_FA2_BA2_IO_021_mb1_FB2_BA2_IO_031,
    input wire        mb1_FA2_BA2_IO_022_mb1_FB2_BA2_IO_008,
    input wire        mb1_FA2_BA2_IO_023_mb1_FB2_BA2_IO_009,
    input wire        mb1_FA2_BA2_IO_024_mb1_FB2_BA2_IO_026,
    input wire        mb1_FA2_BA2_IO_025_mb1_FB2_BA2_IO_027,
    input wire        mb1_FA2_BA2_IO_026_mb1_FB2_BA2_IO_024,
    input wire        mb1_FA2_BA2_IO_027_mb1_FB2_BA2_IO_025,
    input wire        mb1_FA2_BA2_IO_028_mb1_FB2_BA2_IO_042,
    input wire        mb1_FA2_BA2_IO_029_mb1_FB2_BA2_IO_043,
    input wire        mb1_FA2_BA2_IO_030_mb1_FB2_BA2_IO_020,
    input wire        mb1_FA2_BA2_IO_031_mb1_FB2_BA2_IO_021,
    input wire        mb1_FA2_BA2_IO_032_mb1_FB2_BA2_IO_018,
    input wire        mb1_FA2_BA2_IO_033_mb1_FB2_BA2_IO_019,
    input wire        mb1_FA2_BA2_IO_034_mb1_FB2_BA2_IO_036,
    input wire        mb1_FA2_BA2_IO_035_mb1_FB2_BA2_IO_037,
    input wire        mb1_FA2_BA2_IO_036_mb1_FB2_BA2_IO_034,
    input wire        mb1_FA2_BA2_IO_037_mb1_FB2_BA2_IO_035,
    input wire        mb1_FA2_BA2_IO_038_mb1_FB2_BA2_IO_052,
    input wire        mb1_FA2_BA2_IO_039_mb1_FB2_BA2_IO_053,
    input wire        mb1_FA2_BA2_IO_040_mb1_FB2_BA2_IO_050,
    input wire        mb1_FA2_BA2_IO_041_mb1_FB2_BA2_IO_051,
    input wire        mb1_FA2_BA2_IO_042_mb1_FB2_BA2_IO_028,
    input wire        mb1_FA2_BA2_IO_043_mb1_FB2_BA2_IO_029,
    input wire        mb1_FA2_BA2_IO_044_mb1_FB2_BA2_IO_046,
    input wire        mb1_FA2_BA2_IO_045_mb1_FB2_BA2_IO_047,
    input wire        mb1_FA2_BA2_IO_046_mb1_FB2_BA2_IO_044,
    input wire        mb1_FA2_BA2_IO_047_mb1_FB2_BA2_IO_045,
    input wire        mb1_FA2_BA2_IO_048_mb1_FB2_BA2_IO_062,
    input wire        mb1_FA2_BA2_IO_049_mb1_FB2_BA2_IO_063,
    input wire        mb1_FA2_BA2_IO_050_mb1_FB2_BA2_IO_040,
    input wire        mb1_FA2_BA2_IO_051_mb1_FB2_BA2_IO_041,
    input wire        mb1_FA2_BA2_IO_052_mb1_FB2_BA2_IO_038,
    input wire        mb1_FA2_BA2_IO_053_mb1_FB2_BA2_IO_039,
    input wire        mb1_FA2_BA2_IO_054_mb1_FB2_BA2_IO_056,
    input wire        mb1_FA2_BA2_IO_055_mb1_FB2_BA2_IO_057,
    input wire        mb1_FA2_BA2_IO_056_mb1_FB2_BA2_IO_054,
    input wire        mb1_FA2_BA2_IO_057_mb1_FB2_BA2_IO_055,
    input wire        mb1_FA2_BA2_IO_058_mb1_FB2_BA2_IO_072,
    input wire        mb1_FA2_BA2_IO_059_mb1_FB2_BA2_IO_073,
    input wire        mb1_FA2_BA2_IO_060_mb1_FB2_BA2_IO_070,
    input wire        mb1_FA2_BA2_IO_061_mb1_FB2_BA2_IO_071,
    input wire        mb1_FA2_BA2_IO_062_mb1_FB2_BA2_IO_048,
    input wire        mb1_FA2_BA2_IO_063_mb1_FB2_BA2_IO_049,
    input wire        mb1_FA2_BA2_IO_064_mb1_FB2_BA2_IO_066,
    input wire        mb1_FA2_BA2_IO_065_mb1_FB2_BA2_IO_067,
    input wire        mb1_FA2_BA2_IO_066_mb1_FB2_BA2_IO_064,
    input wire        mb1_FA2_BA2_IO_067_mb1_FB2_BA2_IO_065,
    input wire        mb1_FA2_BA2_IO_068_mb1_FB2_BA2_IO_082,
    input wire        mb1_FA2_BA2_IO_069_mb1_FB2_BA2_IO_083,
    input wire        mb1_FA2_BA2_IO_070_mb1_FB2_BA2_IO_060,
    input wire        mb1_FA2_BA2_IO_071_mb1_FB2_BA2_IO_061,
    input wire        mb1_FA2_BA2_IO_072_mb1_FB2_BA2_IO_058,
    input wire        mb1_FA2_BA2_IO_073_mb1_FB2_BA2_IO_059,
    input wire        mb1_FA2_BA2_IO_074_mb1_FB2_BA2_IO_076,
    input wire        mb1_FA2_BA2_IO_075_mb1_FB2_BA2_IO_077,
    input wire        mb1_FA2_BA2_IO_076_mb1_FB2_BA2_IO_074,
    input wire        mb1_FA2_BA2_IO_077_mb1_FB2_BA2_IO_075,
    input wire        mb1_FA2_BA2_IO_078_mb1_FB2_BA2_IO_092,
    input wire        mb1_FA2_BA2_IO_079_mb1_FB2_BA2_IO_093,
    input wire        mb1_FA2_BA2_IO_080_mb1_FB2_BA2_IO_090,
    input wire        mb1_FA2_BA2_IO_081_mb1_FB2_BA2_IO_091,
    input wire        mb1_FA2_BA2_IO_082_mb1_FB2_BA2_IO_068,
    input wire        mb1_FA2_BA2_IO_083_mb1_FB2_BA2_IO_069,
    input wire        mb1_FA2_BA2_IO_084_mb1_FB2_BA2_IO_086,
    input wire        mb1_FA2_BA2_IO_085_mb1_FB2_BA2_IO_087,
    input wire        mb1_FA2_BA2_IO_086_mb1_FB2_BA2_IO_084,
    input wire        mb1_FA2_BA2_IO_087_mb1_FB2_BA2_IO_085,
    input wire        mb1_FA2_BA2_IO_088_mb1_FB2_BA2_IO_102,
    input wire        mb1_FA2_BA2_IO_089_mb1_FB2_BA2_IO_103,
    input wire        mb1_FA2_BA2_IO_090_mb1_FB2_BA2_IO_080,
    input wire        mb1_FA2_BA2_IO_091_mb1_FB2_BA2_IO_081,
    input wire        mb1_FA2_BA2_IO_092_mb1_FB2_BA2_IO_078,
    input wire        mb1_FA2_BA2_IO_093_mb1_FB2_BA2_IO_079,
    input wire        mb1_FA2_BA2_IO_094_mb1_FB2_BA2_IO_096,
    input wire        mb1_FA2_BA2_IO_095_mb1_FB2_BA2_IO_097,
    input wire        mb1_FA2_BA2_IO_096_mb1_FB2_BA2_IO_094,
    input wire        mb1_FA2_BA2_IO_097_mb1_FB2_BA2_IO_095,
    input wire        mb1_FA2_BA2_IO_098_mb1_FB2_BA2_IO_112,
    input wire        mb1_FA2_BA2_IO_099_mb1_FB2_BA2_IO_113,
    input wire        mb1_FA2_BA2_IO_100_mb1_FB2_BA2_IO_110,
    input wire        mb1_FA2_BA2_IO_101_mb1_FB2_BA2_IO_111,
    input wire        mb1_FA2_BA2_IO_102_mb1_FB2_BA2_IO_088,
    input wire        mb1_FA2_BA2_IO_103_mb1_FB2_BA2_IO_089,
    input wire        mb1_FA2_BA2_IO_104_mb1_FB2_BA2_IO_106,
    input wire        mb1_FA2_BA2_IO_105_mb1_FB2_BA2_IO_107,
    input wire        mb1_FA2_BA2_IO_106_mb1_FB2_BA2_IO_104,
    input wire        mb1_FA2_BA2_IO_107_mb1_FB2_BA2_IO_105,
    input wire        mb1_FA2_BA2_IO_108_mb1_FB2_BA2_IO_122,
    input wire        mb1_FA2_BA2_IO_109_mb1_FB2_BA2_IO_123,
    input wire        mb1_FA2_BA2_IO_110_mb1_FB2_BA2_IO_100,
    input wire        mb1_FA2_BA2_IO_111_mb1_FB2_BA2_IO_101,
    input wire        mb1_FA2_BA2_IO_112_mb1_FB2_BA2_IO_098,
    input wire        mb1_FA2_BA2_IO_113_mb1_FB2_BA2_IO_099,
    input wire        mb1_FA2_BA2_IO_114_mb1_FB2_BA2_IO_116,
    input wire        mb1_FA2_BA2_IO_115_mb1_FB2_BA2_IO_117,
    input wire        mb1_FA2_BA2_IO_116_mb1_FB2_BA2_IO_114,
    input wire        mb1_FA2_BA2_IO_117_mb1_FB2_BA2_IO_115,
    input wire        mb1_FA2_BA2_IO_118_mb1_FB2_BA2_IO_132,
    input wire        mb1_FA2_BA2_IO_119_mb1_FB2_BA2_IO_133,
    input wire        mb1_FA2_BA2_IO_120_mb1_FB2_BA2_IO_130,
    input wire        mb1_FA2_BA2_IO_121_mb1_FB2_BA2_IO_131,
    input wire        mb1_FA2_BA2_IO_122_mb1_FB2_BA2_IO_108,
    input wire        mb1_FA2_BA2_IO_123_mb1_FB2_BA2_IO_109,
    input wire        mb1_FA2_BA2_IO_124_mb1_FB2_BA2_IO_126,
    input wire        mb1_FA2_BA2_IO_125_mb1_FB2_BA2_IO_127,
    input wire        mb1_FA2_BA2_IO_126_mb1_FB2_BA2_IO_124,
    input wire        mb1_FA2_BA2_IO_127_mb1_FB2_BA2_IO_125,
    input wire        mb1_FA2_BA2_IO_130_mb1_FB2_BA2_IO_120,
    input wire        mb1_FA2_BA2_IO_131_mb1_FB2_BA2_IO_121,
    input wire        mb1_FA2_BA2_IO_132_mb1_FB2_BA2_IO_118,
    input wire        mb1_FA2_BA2_IO_133_mb1_FB2_BA2_IO_119,
    input wire        mb1_FA2_BA2_IO_134_mb1_FB2_BA2_IO_136,
    input wire        mb1_FA2_BA2_IO_136_mb1_FB2_BA2_IO_134,
    input wire        mb1_FB1_TA1_CLKIO_N_0_mb1_FB2_BB0_CLKIO_N_7,
    input wire        mb1_FB1_TA1_CLKIO_N_1_mb1_FB2_BB0_CLKIO_N_6,
    input wire        mb1_FB1_TA1_CLKIO_N_2_mb1_FB2_BB0_CLKIO_N_4,
    input wire        mb1_FB1_TA1_CLKIO_N_3_mb1_FB2_BB0_CLKIO_N_3,
    input wire        mb1_FB1_TA1_CLKIO_N_4_mb1_FB2_BB0_CLKIO_N_2,
    input wire        mb1_FB1_TA1_CLKIO_N_5_mb1_FB2_BB0_IO_010,
    input wire        mb1_FB1_TA1_CLKIO_N_6_mb1_FB2_BB0_CLKIO_N_1,
    input wire        mb1_FB1_TA1_CLKIO_N_7_mb1_FB2_BB0_CLKIO_N_0,
    input wire        mb1_FB1_TA1_CLKIO_P_0_mb1_FB2_BB0_CLKIO_P_7,
    input wire        mb1_FB1_TA1_CLKIO_P_1_mb1_FB2_BB0_CLKIO_P_6,
    input wire        mb1_FB1_TA1_CLKIO_P_2_mb1_FB2_BB0_CLKIO_P_4,
    input wire        mb1_FB1_TA1_CLKIO_P_3_mb1_FB2_BB0_CLKIO_P_3,
    input wire        mb1_FB1_TA1_CLKIO_P_4_mb1_FB2_BB0_CLKIO_P_2,
    input wire        mb1_FB1_TA1_CLKIO_P_5_mb1_FB2_BB0_IO_011,
    input wire        mb1_FB1_TA1_CLKIO_P_6_mb1_FB2_BB0_CLKIO_P_1,
    input wire        mb1_FB1_TA1_CLKIO_P_7_mb1_FB2_BB0_CLKIO_P_0,
    input wire        mb1_FB1_TA1_IO_004_mb1_FB2_BB0_IO_006,
    input wire        mb1_FB1_TA1_IO_005_mb1_FB2_BB0_IO_007,
    input wire        mb1_FB1_TA1_IO_006_mb1_FB2_BB0_IO_004,
    input wire        mb1_FB1_TA1_IO_007_mb1_FB2_BB0_IO_005,
    input wire        mb1_FB1_TA1_IO_008_mb1_FB2_BB0_IO_022,
    input wire        mb1_FB1_TA1_IO_009_mb1_FB2_BB0_IO_023,
    input wire        mb1_FB1_TA1_IO_010_mb1_FB2_BB0_CLKIO_N_5,
    input wire        mb1_FB1_TA1_IO_011_mb1_FB2_BB0_CLKIO_P_5,
    input wire        mb1_FB1_TA1_IO_012_mb1_FB2_BB0_IO_012,
    input wire        mb1_FB1_TA1_IO_013_mb1_FB2_BB0_IO_013,
    input wire        mb1_FB1_TA1_IO_014_mb1_FB2_BB0_IO_016,
    input wire        mb1_FB1_TA1_IO_015_mb1_FB2_BB0_IO_017,
    input wire        mb1_FB1_TA1_IO_016_mb1_FB2_BB0_IO_014,
    input wire        mb1_FB1_TA1_IO_017_mb1_FB2_BB0_IO_015,
    input wire        mb1_FB1_TA1_IO_018_mb1_FB2_BB0_IO_032,
    input wire        mb1_FB1_TA1_IO_019_mb1_FB2_BB0_IO_033,
    input wire        mb1_FB1_TA1_IO_020_mb1_FB2_BB0_IO_030,
    input wire        mb1_FB1_TA1_IO_021_mb1_FB2_BB0_IO_031,
    input wire        mb1_FB1_TA1_IO_022_mb1_FB2_BB0_IO_008,
    input wire        mb1_FB1_TA1_IO_023_mb1_FB2_BB0_IO_009,
    input wire        mb1_FB1_TA1_IO_024_mb1_FB2_BB0_IO_026,
    input wire        mb1_FB1_TA1_IO_025_mb1_FB2_BB0_IO_027,
    input wire        mb1_FB1_TA1_IO_026_mb1_FB2_BB0_IO_024,
    input wire        mb1_FB1_TA1_IO_027_mb1_FB2_BB0_IO_025,
    input wire        mb1_FB1_TA1_IO_028_mb1_FB2_BB0_IO_042,
    input wire        mb1_FB1_TA1_IO_029_mb1_FB2_BB0_IO_043,
    input wire        mb1_FB1_TA1_IO_030_mb1_FB2_BB0_IO_020,
    input wire        mb1_FB1_TA1_IO_031_mb1_FB2_BB0_IO_021,
    input wire        mb1_FB1_TA1_IO_032_mb1_FB2_BB0_IO_018,
    input wire        mb1_FB1_TA1_IO_033_mb1_FB2_BB0_IO_019,
    input wire        mb1_FB1_TA1_IO_034_mb1_FB2_BB0_IO_036,
    input wire        mb1_FB1_TA1_IO_035_mb1_FB2_BB0_IO_037,
    input wire        mb1_FB1_TA1_IO_036_mb1_FB2_BB0_IO_034,
    input wire        mb1_FB1_TA1_IO_037_mb1_FB2_BB0_IO_035,
    input wire        mb1_FB1_TA1_IO_038_mb1_FB2_BB0_IO_052,
    input wire        mb1_FB1_TA1_IO_039_mb1_FB2_BB0_IO_053,
    input wire        mb1_FB1_TA1_IO_040_mb1_FB2_BB0_IO_050,
    input wire        mb1_FB1_TA1_IO_041_mb1_FB2_BB0_IO_051,
    input wire        mb1_FB1_TA1_IO_042_mb1_FB2_BB0_IO_028,
    input wire        mb1_FB1_TA1_IO_043_mb1_FB2_BB0_IO_029,
    input wire        mb1_FB1_TA1_IO_044_mb1_FB2_BB0_IO_046,
    input wire        mb1_FB1_TA1_IO_045_mb1_FB2_BB0_IO_047,
    input wire        mb1_FB1_TA1_IO_046_mb1_FB2_BB0_IO_044,
    input wire        mb1_FB1_TA1_IO_047_mb1_FB2_BB0_IO_045,
    input wire        mb1_FB1_TA1_IO_048_mb1_FB2_BB0_IO_062,
    input wire        mb1_FB1_TA1_IO_049_mb1_FB2_BB0_IO_063,
    input wire        mb1_FB1_TA1_IO_050_mb1_FB2_BB0_IO_040,
    input wire        mb1_FB1_TA1_IO_051_mb1_FB2_BB0_IO_041,
    input wire        mb1_FB1_TA1_IO_052_mb1_FB2_BB0_IO_038,
    input wire        mb1_FB1_TA1_IO_053_mb1_FB2_BB0_IO_039,
    input wire        mb1_FB1_TA1_IO_054_mb1_FB2_BB0_IO_056,
    input wire        mb1_FB1_TA1_IO_055_mb1_FB2_BB0_IO_057,
    input wire        mb1_FB1_TA1_IO_056_mb1_FB2_BB0_IO_054,
    input wire        mb1_FB1_TA1_IO_057_mb1_FB2_BB0_IO_055,
    input wire        mb1_FB1_TA1_IO_058_mb1_FB2_BB0_IO_072,
    input wire        mb1_FB1_TA1_IO_059_mb1_FB2_BB0_IO_073,
    input wire        mb1_FB1_TA1_IO_060_mb1_FB2_BB0_IO_070,
    input wire        mb1_FB1_TA1_IO_061_mb1_FB2_BB0_IO_071,
    input wire        mb1_FB1_TA1_IO_062_mb1_FB2_BB0_IO_048,
    input wire        mb1_FB1_TA1_IO_063_mb1_FB2_BB0_IO_049,
    input wire        mb1_FB1_TA1_IO_064_mb1_FB2_BB0_IO_066,
    input wire        mb1_FB1_TA1_IO_065_mb1_FB2_BB0_IO_067,
    input wire        mb1_FB1_TA1_IO_066_mb1_FB2_BB0_IO_064,
    input wire        mb1_FB1_TA1_IO_067_mb1_FB2_BB0_IO_065,
    input wire        mb1_FB1_TA1_IO_068_mb1_FB2_BB0_IO_082,
    input wire        mb1_FB1_TA1_IO_069_mb1_FB2_BB0_IO_083,
    input wire        mb1_FB1_TA1_IO_070_mb1_FB2_BB0_IO_060,
    input wire        mb1_FB1_TA1_IO_071_mb1_FB2_BB0_IO_061,
    input wire        mb1_FB1_TA1_IO_072_mb1_FB2_BB0_IO_058,
    input wire        mb1_FB1_TA1_IO_073_mb1_FB2_BB0_IO_059,
    input wire        mb1_FB1_TA1_IO_074_mb1_FB2_BB0_IO_076,
    input wire        mb1_FB1_TA1_IO_075_mb1_FB2_BB0_IO_077,
    input wire        mb1_FB1_TA1_IO_076_mb1_FB2_BB0_IO_074,
    input wire        mb1_FB1_TA1_IO_077_mb1_FB2_BB0_IO_075,
    input wire        mb1_FB1_TA1_IO_078_mb1_FB2_BB0_IO_092,
    input wire        mb1_FB1_TA1_IO_079_mb1_FB2_BB0_IO_093,
    input wire        mb1_FB1_TA1_IO_080_mb1_FB2_BB0_IO_090,
    input wire        mb1_FB1_TA1_IO_081_mb1_FB2_BB0_IO_091,
    input wire        mb1_FB1_TA1_IO_082_mb1_FB2_BB0_IO_068,
    input wire        mb1_FB1_TA1_IO_083_mb1_FB2_BB0_IO_069,
    input wire        mb1_FB1_TA1_IO_084_mb1_FB2_BB0_IO_086,
    input wire        mb1_FB1_TA1_IO_085_mb1_FB2_BB0_IO_087,
    input wire        mb1_FB1_TA1_IO_086_mb1_FB2_BB0_IO_084,
    input wire        mb1_FB1_TA1_IO_087_mb1_FB2_BB0_IO_085,
    input wire        mb1_FB1_TA1_IO_088_mb1_FB2_BB0_IO_102,
    input wire        mb1_FB1_TA1_IO_089_mb1_FB2_BB0_IO_103,
    input wire        mb1_FB1_TA1_IO_090_mb1_FB2_BB0_IO_080,
    input wire        mb1_FB1_TA1_IO_091_mb1_FB2_BB0_IO_081,
    input wire        mb1_FB1_TA1_IO_092_mb1_FB2_BB0_IO_078,
    input wire        mb1_FB1_TA1_IO_093_mb1_FB2_BB0_IO_079,
    input wire        mb1_FB1_TA1_IO_094_mb1_FB2_BB0_IO_096,
    input wire        mb1_FB1_TA1_IO_095_mb1_FB2_BB0_IO_097,
    input wire        mb1_FB1_TA1_IO_096_mb1_FB2_BB0_IO_094,
    input wire        mb1_FB1_TA1_IO_097_mb1_FB2_BB0_IO_095,
    input wire        mb1_FB1_TA1_IO_098_mb1_FB2_BB0_IO_112,
    input wire        mb1_FB1_TA1_IO_099_mb1_FB2_BB0_IO_113,
    input wire        mb1_FB1_TA1_IO_100_mb1_FB2_BB0_IO_110,
    input wire        mb1_FB1_TA1_IO_101_mb1_FB2_BB0_IO_111,
    input wire        mb1_FB1_TA1_IO_102_mb1_FB2_BB0_IO_088,
    input wire        mb1_FB1_TA1_IO_103_mb1_FB2_BB0_IO_089,
    input wire        mb1_FB1_TA1_IO_104_mb1_FB2_BB0_IO_106,
    input wire        mb1_FB1_TA1_IO_105_mb1_FB2_BB0_IO_107,
    input wire        mb1_FB1_TA1_IO_106_mb1_FB2_BB0_IO_104,
    input wire        mb1_FB1_TA1_IO_107_mb1_FB2_BB0_IO_105,
    input wire        mb1_FB1_TA1_IO_108_mb1_FB2_BB0_IO_122,
    input wire        mb1_FB1_TA1_IO_109_mb1_FB2_BB0_IO_123,
    input wire        mb1_FB1_TA1_IO_110_mb1_FB2_BB0_IO_100,
    input wire        mb1_FB1_TA1_IO_111_mb1_FB2_BB0_IO_101,
    input wire        mb1_FB1_TA1_IO_112_mb1_FB2_BB0_IO_098,
    input wire        mb1_FB1_TA1_IO_113_mb1_FB2_BB0_IO_099,
    input wire        mb1_FB1_TA1_IO_114_mb1_FB2_BB0_IO_116,
    input wire        mb1_FB1_TA1_IO_115_mb1_FB2_BB0_IO_117,
    input wire        mb1_FB1_TA1_IO_116_mb1_FB2_BB0_IO_114,
    input wire        mb1_FB1_TA1_IO_117_mb1_FB2_BB0_IO_115,
    input wire        mb1_FB1_TA1_IO_118_mb1_FB2_BB0_IO_132,
    input wire        mb1_FB1_TA1_IO_119_mb1_FB2_BB0_IO_133,
    input wire        mb1_FB1_TA1_IO_120_mb1_FB2_BB0_IO_130,
    input wire        mb1_FB1_TA1_IO_121_mb1_FB2_BB0_IO_131,
    input wire        mb1_FB1_TA1_IO_122_mb1_FB2_BB0_IO_108,
    input wire        mb1_FB1_TA1_IO_123_mb1_FB2_BB0_IO_109,
    input wire        mb1_FB1_TA1_IO_124_mb1_FB2_BB0_IO_126,
    input wire        mb1_FB1_TA1_IO_125_mb1_FB2_BB0_IO_127,
    input wire        mb1_FB1_TA1_IO_126_mb1_FB2_BB0_IO_124,
    input wire        mb1_FB1_TA1_IO_127_mb1_FB2_BB0_IO_125,
    input wire        mb1_FB1_TA1_IO_130_mb1_FB2_BB0_IO_120,
    input wire        mb1_FB1_TA1_IO_131_mb1_FB2_BB0_IO_121,
    input wire        mb1_FB1_TA1_IO_132_mb1_FB2_BB0_IO_118,
    input wire        mb1_FB1_TA1_IO_133_mb1_FB2_BB0_IO_119,
    input wire        mb1_FB1_TA1_IO_134_mb1_FB2_BB0_IO_136,
    input wire        mb1_FB1_TA1_IO_136_mb1_FB2_BB0_IO_134,
    input wire        mb1_FA1_TB2_CLKIO_N_0_mb1_FB2_BB1_CLKIO_N_7,
    input wire        mb1_FA1_TB2_CLKIO_N_1_mb1_FB2_BB1_CLKIO_N_6,
    input wire        mb1_FA1_TB2_CLKIO_N_2_mb1_FB2_BB1_CLKIO_N_4,
    input wire        mb1_FA1_TB2_CLKIO_N_3_mb1_FB2_BB1_CLKIO_N_3,
    input wire        mb1_FA1_TB2_CLKIO_N_4_mb1_FB2_BB1_CLKIO_N_2,
    input wire        mb1_FA1_TB2_CLKIO_N_5_mb1_FB2_BB1_IO_010,
    input wire        mb1_FA1_TB2_CLKIO_N_6_mb1_FB2_BB1_CLKIO_N_1,
    input wire        mb1_FA1_TB2_CLKIO_N_7_mb1_FB2_BB1_CLKIO_N_0,
    input wire        mb1_FA1_TB2_CLKIO_P_0_mb1_FB2_BB1_CLKIO_P_7,
    input wire        mb1_FA1_TB2_CLKIO_P_1_mb1_FB2_BB1_CLKIO_P_6,
    input wire        mb1_FA1_TB2_CLKIO_P_2_mb1_FB2_BB1_CLKIO_P_4,
    input wire        mb1_FA1_TB2_CLKIO_P_3_mb1_FB2_BB1_CLKIO_P_3,
    input wire        mb1_FA1_TB2_CLKIO_P_4_mb1_FB2_BB1_CLKIO_P_2,
    input wire        mb1_FA1_TB2_CLKIO_P_5_mb1_FB2_BB1_IO_011,
    input wire        mb1_FA1_TB2_CLKIO_P_6_mb1_FB2_BB1_CLKIO_P_1,
    input wire        mb1_FA1_TB2_CLKIO_P_7_mb1_FB2_BB1_CLKIO_P_0,
    input wire        mb1_FA1_TB2_IO_004_mb1_FB2_BB1_IO_006,
    input wire        mb1_FA1_TB2_IO_005_mb1_FB2_BB1_IO_007,
    input wire        mb1_FA1_TB2_IO_006_mb1_FB2_BB1_IO_004,
    input wire        mb1_FA1_TB2_IO_007_mb1_FB2_BB1_IO_005,
    input wire        mb1_FA1_TB2_IO_008_mb1_FB2_BB1_IO_022,
    input wire        mb1_FA1_TB2_IO_009_mb1_FB2_BB1_IO_023,
    input wire        mb1_FA1_TB2_IO_010_mb1_FB2_BB1_CLKIO_N_5,
    input wire        mb1_FA1_TB2_IO_011_mb1_FB2_BB1_CLKIO_P_5,
    input wire        mb1_FA1_TB2_IO_012_mb1_FB2_BB1_IO_012,
    input wire        mb1_FA1_TB2_IO_013_mb1_FB2_BB1_IO_013,
    input wire        mb1_FA1_TB2_IO_014_mb1_FB2_BB1_IO_016,
    input wire        mb1_FA1_TB2_IO_015_mb1_FB2_BB1_IO_017,
    input wire        mb1_FA1_TB2_IO_016_mb1_FB2_BB1_IO_014,
    input wire        mb1_FA1_TB2_IO_017_mb1_FB2_BB1_IO_015,
    input wire        mb1_FA1_TB2_IO_018_mb1_FB2_BB1_IO_032,
    input wire        mb1_FA1_TB2_IO_019_mb1_FB2_BB1_IO_033,
    input wire        mb1_FA1_TB2_IO_020_mb1_FB2_BB1_IO_030,
    input wire        mb1_FA1_TB2_IO_021_mb1_FB2_BB1_IO_031,
    input wire        mb1_FA1_TB2_IO_022_mb1_FB2_BB1_IO_008,
    input wire        mb1_FA1_TB2_IO_023_mb1_FB2_BB1_IO_009,
    input wire        mb1_FA1_TB2_IO_024_mb1_FB2_BB1_IO_026,
    input wire        mb1_FA1_TB2_IO_025_mb1_FB2_BB1_IO_027,
    input wire        mb1_FA1_TB2_IO_026_mb1_FB2_BB1_IO_024,
    input wire        mb1_FA1_TB2_IO_027_mb1_FB2_BB1_IO_025,
    input wire        mb1_FA1_TB2_IO_028_mb1_FB2_BB1_IO_042,
    input wire        mb1_FA1_TB2_IO_029_mb1_FB2_BB1_IO_043,
    input wire        mb1_FA1_TB2_IO_030_mb1_FB2_BB1_IO_020,
    input wire        mb1_FA1_TB2_IO_031_mb1_FB2_BB1_IO_021,
    input wire        mb1_FA1_TB2_IO_032_mb1_FB2_BB1_IO_018,
    input wire        mb1_FA1_TB2_IO_033_mb1_FB2_BB1_IO_019,
    input wire        mb1_FA1_TB2_IO_034_mb1_FB2_BB1_IO_036,
    input wire        mb1_FA1_TB2_IO_035_mb1_FB2_BB1_IO_037,
    input wire        mb1_FA1_TB2_IO_036_mb1_FB2_BB1_IO_034,
    input wire        mb1_FA1_TB2_IO_037_mb1_FB2_BB1_IO_035,
    input wire        mb1_FA1_TB2_IO_038_mb1_FB2_BB1_IO_052,
    input wire        mb1_FA1_TB2_IO_039_mb1_FB2_BB1_IO_053,
    input wire        mb1_FA1_TB2_IO_040_mb1_FB2_BB1_IO_050,
    input wire        mb1_FA1_TB2_IO_041_mb1_FB2_BB1_IO_051,
    input wire        mb1_FA1_TB2_IO_042_mb1_FB2_BB1_IO_028,
    input wire        mb1_FA1_TB2_IO_043_mb1_FB2_BB1_IO_029,
    input wire        mb1_FA1_TB2_IO_044_mb1_FB2_BB1_IO_046,
    input wire        mb1_FA1_TB2_IO_045_mb1_FB2_BB1_IO_047,
    input wire        mb1_FA1_TB2_IO_046_mb1_FB2_BB1_IO_044,
    input wire        mb1_FA1_TB2_IO_047_mb1_FB2_BB1_IO_045,
    input wire        mb1_FA1_TB2_IO_048_mb1_FB2_BB1_IO_062,
    input wire        mb1_FA1_TB2_IO_049_mb1_FB2_BB1_IO_063,
    input wire        mb1_FA1_TB2_IO_050_mb1_FB2_BB1_IO_040,
    input wire        mb1_FA1_TB2_IO_051_mb1_FB2_BB1_IO_041,
    input wire        mb1_FA1_TB2_IO_052_mb1_FB2_BB1_IO_038,
    input wire        mb1_FA1_TB2_IO_053_mb1_FB2_BB1_IO_039,
    input wire        mb1_FA1_TB2_IO_054_mb1_FB2_BB1_IO_056,
    input wire        mb1_FA1_TB2_IO_055_mb1_FB2_BB1_IO_057,
    input wire        mb1_FA1_TB2_IO_056_mb1_FB2_BB1_IO_054,
    input wire        mb1_FA1_TB2_IO_057_mb1_FB2_BB1_IO_055,
    input wire        mb1_FA1_TB2_IO_058_mb1_FB2_BB1_IO_072,
    input wire        mb1_FA1_TB2_IO_059_mb1_FB2_BB1_IO_073,
    input wire        mb1_FA1_TB2_IO_060_mb1_FB2_BB1_IO_070,
    input wire        mb1_FA1_TB2_IO_061_mb1_FB2_BB1_IO_071,
    input wire        mb1_FA1_TB2_IO_062_mb1_FB2_BB1_IO_048,
    input wire        mb1_FA1_TB2_IO_063_mb1_FB2_BB1_IO_049,
    input wire        mb1_FA1_TB2_IO_064_mb1_FB2_BB1_IO_066,
    input wire        mb1_FA1_TB2_IO_065_mb1_FB2_BB1_IO_067,
    input wire        mb1_FA1_TB2_IO_066_mb1_FB2_BB1_IO_064,
    input wire        mb1_FA1_TB2_IO_067_mb1_FB2_BB1_IO_065,
    input wire        mb1_FA1_TB2_IO_068_mb1_FB2_BB1_IO_082,
    input wire        mb1_FA1_TB2_IO_069_mb1_FB2_BB1_IO_083,
    input wire        mb1_FA1_TB2_IO_070_mb1_FB2_BB1_IO_060,
    input wire        mb1_FA1_TB2_IO_071_mb1_FB2_BB1_IO_061,
    input wire        mb1_FA1_TB2_IO_072_mb1_FB2_BB1_IO_058,
    input wire        mb1_FA1_TB2_IO_073_mb1_FB2_BB1_IO_059,
    input wire        mb1_FA1_TB2_IO_074_mb1_FB2_BB1_IO_076,
    input wire        mb1_FA1_TB2_IO_075_mb1_FB2_BB1_IO_077,
    input wire        mb1_FA1_TB2_IO_076_mb1_FB2_BB1_IO_074,
    input wire        mb1_FA1_TB2_IO_077_mb1_FB2_BB1_IO_075,
    input wire        mb1_FA1_TB2_IO_078_mb1_FB2_BB1_IO_092,
    input wire        mb1_FA1_TB2_IO_079_mb1_FB2_BB1_IO_093,
    input wire        mb1_FA1_TB2_IO_080_mb1_FB2_BB1_IO_090,
    input wire        mb1_FA1_TB2_IO_081_mb1_FB2_BB1_IO_091,
    input wire        mb1_FA1_TB2_IO_082_mb1_FB2_BB1_IO_068,
    input wire        mb1_FA1_TB2_IO_083_mb1_FB2_BB1_IO_069,
    input wire        mb1_FA1_TB2_IO_084_mb1_FB2_BB1_IO_086,
    input wire        mb1_FA1_TB2_IO_085_mb1_FB2_BB1_IO_087,
    input wire        mb1_FA1_TB2_IO_086_mb1_FB2_BB1_IO_084,
    input wire        mb1_FA1_TB2_IO_087_mb1_FB2_BB1_IO_085,
    input wire        mb1_FA1_TB2_IO_088_mb1_FB2_BB1_IO_102,
    input wire        mb1_FA1_TB2_IO_089_mb1_FB2_BB1_IO_103,
    input wire        mb1_FA1_TB2_IO_090_mb1_FB2_BB1_IO_080,
    input wire        mb1_FA1_TB2_IO_091_mb1_FB2_BB1_IO_081,
    input wire        mb1_FA1_TB2_IO_092_mb1_FB2_BB1_IO_078,
    input wire        mb1_FA1_TB2_IO_093_mb1_FB2_BB1_IO_079,
    input wire        mb1_FA1_TB2_IO_094_mb1_FB2_BB1_IO_096,
    input wire        mb1_FA1_TB2_IO_095_mb1_FB2_BB1_IO_097,
    input wire        mb1_FA1_TB2_IO_096_mb1_FB2_BB1_IO_094,
    input wire        mb1_FA1_TB2_IO_097_mb1_FB2_BB1_IO_095,
    input wire        mb1_FA1_TB2_IO_098_mb1_FB2_BB1_IO_112,
    input wire        mb1_FA1_TB2_IO_099_mb1_FB2_BB1_IO_113,
    input wire        mb1_FA1_TB2_IO_100_mb1_FB2_BB1_IO_110,
    input wire        mb1_FA1_TB2_IO_101_mb1_FB2_BB1_IO_111,
    input wire        mb1_FA1_TB2_IO_102_mb1_FB2_BB1_IO_088,
    input wire        mb1_FA1_TB2_IO_103_mb1_FB2_BB1_IO_089,
    input wire        mb1_FA1_TB2_IO_104_mb1_FB2_BB1_IO_106,
    input wire        mb1_FA1_TB2_IO_105_mb1_FB2_BB1_IO_107,
    input wire        mb1_FA1_TB2_IO_106_mb1_FB2_BB1_IO_104,
    input wire        mb1_FA1_TB2_IO_107_mb1_FB2_BB1_IO_105,
    input wire        mb1_FA1_TB2_IO_108_mb1_FB2_BB1_IO_122,
    input wire        mb1_FA1_TB2_IO_109_mb1_FB2_BB1_IO_123,
    input wire        mb1_FA1_TB2_IO_110_mb1_FB2_BB1_IO_100,
    input wire        mb1_FA1_TB2_IO_111_mb1_FB2_BB1_IO_101,
    input wire        mb1_FA1_TB2_IO_112_mb1_FB2_BB1_IO_098,
    input wire        mb1_FA1_TB2_IO_113_mb1_FB2_BB1_IO_099,
    input wire        mb1_FA1_TB2_IO_114_mb1_FB2_BB1_IO_116,
    input wire        mb1_FA1_TB2_IO_115_mb1_FB2_BB1_IO_117,
    input wire        mb1_FA1_TB2_IO_116_mb1_FB2_BB1_IO_114,
    input wire        mb1_FA1_TB2_IO_117_mb1_FB2_BB1_IO_115,
    input wire        mb1_FA1_TB2_IO_118_mb1_FB2_BB1_IO_132,
    input wire        mb1_FA1_TB2_IO_119_mb1_FB2_BB1_IO_133,
    input wire        mb1_FA1_TB2_IO_120_mb1_FB2_BB1_IO_130,
    input wire        mb1_FA1_TB2_IO_121_mb1_FB2_BB1_IO_131,
    input wire        mb1_FA1_TB2_IO_122_mb1_FB2_BB1_IO_108,
    input wire        mb1_FA1_TB2_IO_123_mb1_FB2_BB1_IO_109,
    input wire        mb1_FA1_TB2_IO_124_mb1_FB2_BB1_IO_126,
    input wire        mb1_FA1_TB2_IO_125_mb1_FB2_BB1_IO_127,
    input wire        mb1_FA1_TB2_IO_126_mb1_FB2_BB1_IO_124,
    input wire        mb1_FA1_TB2_IO_127_mb1_FB2_BB1_IO_125,
    input wire        mb1_FA1_TB2_IO_130_mb1_FB2_BB1_IO_120,
    input wire        mb1_FA1_TB2_IO_131_mb1_FB2_BB1_IO_121,
    input wire        mb1_FA1_TB2_IO_132_mb1_FB2_BB1_IO_118,
    input wire        mb1_FA1_TB2_IO_133_mb1_FB2_BB1_IO_119,
    input wire        mb1_FA1_TB2_IO_134_mb1_FB2_BB1_IO_136,
    input wire        mb1_FA1_TB2_IO_136_mb1_FB2_BB1_IO_134,
    input wire        mb1_FB1_TB0_CLKIO_N_0_mb1_FB2_BB2_CLKIO_N_7,
    input wire        mb1_FB1_TB0_CLKIO_N_1_mb1_FB2_BB2_CLKIO_N_6,
    input wire        mb1_FB1_TB0_CLKIO_N_2_mb1_FB2_BB2_CLKIO_N_4,
    input wire        mb1_FB1_TB0_CLKIO_N_3_mb1_FB2_BB2_CLKIO_N_3,
    input wire        mb1_FB1_TB0_CLKIO_N_4_mb1_FB2_BB2_CLKIO_N_2,
    input wire        mb1_FB1_TB0_CLKIO_N_5_mb1_FB2_BB2_IO_010,
    input wire        mb1_FB1_TB0_CLKIO_N_6_mb1_FB2_BB2_CLKIO_N_1,
    input wire        mb1_FB1_TB0_CLKIO_N_7_mb1_FB2_BB2_CLKIO_N_0,
    input wire        mb1_FB1_TB0_CLKIO_P_0_mb1_FB2_BB2_CLKIO_P_7,
    input wire        mb1_FB1_TB0_CLKIO_P_1_mb1_FB2_BB2_CLKIO_P_6,
    input wire        mb1_FB1_TB0_CLKIO_P_2_mb1_FB2_BB2_CLKIO_P_4,
    input wire        mb1_FB1_TB0_CLKIO_P_3_mb1_FB2_BB2_CLKIO_P_3,
    input wire        mb1_FB1_TB0_CLKIO_P_4_mb1_FB2_BB2_CLKIO_P_2,
    input wire        mb1_FB1_TB0_CLKIO_P_5_mb1_FB2_BB2_IO_011,
    input wire        mb1_FB1_TB0_CLKIO_P_6_mb1_FB2_BB2_CLKIO_P_1,
    input wire        mb1_FB1_TB0_CLKIO_P_7_mb1_FB2_BB2_CLKIO_P_0,
    input wire        mb1_FB1_TB0_IO_004_mb1_FB2_BB2_IO_006,
    input wire        mb1_FB1_TB0_IO_005_mb1_FB2_BB2_IO_007,
    input wire        mb1_FB1_TB0_IO_006_mb1_FB2_BB2_IO_004,
    input wire        mb1_FB1_TB0_IO_007_mb1_FB2_BB2_IO_005,
    input wire        mb1_FB1_TB0_IO_008_mb1_FB2_BB2_IO_022,
    input wire        mb1_FB1_TB0_IO_009_mb1_FB2_BB2_IO_023,
    input wire        mb1_FB1_TB0_IO_010_mb1_FB2_BB2_CLKIO_N_5,
    input wire        mb1_FB1_TB0_IO_011_mb1_FB2_BB2_CLKIO_P_5,
    input wire        mb1_FB1_TB0_IO_012_mb1_FB2_BB2_IO_012,
    input wire        mb1_FB1_TB0_IO_013_mb1_FB2_BB2_IO_013,
    input wire        mb1_FB1_TB0_IO_014_mb1_FB2_BB2_IO_016,
    input wire        mb1_FB1_TB0_IO_015_mb1_FB2_BB2_IO_017,
    input wire        mb1_FB1_TB0_IO_016_mb1_FB2_BB2_IO_014,
    input wire        mb1_FB1_TB0_IO_017_mb1_FB2_BB2_IO_015,
    input wire        mb1_FB1_TB0_IO_018_mb1_FB2_BB2_IO_032,
    input wire        mb1_FB1_TB0_IO_019_mb1_FB2_BB2_IO_033,
    input wire        mb1_FB1_TB0_IO_020_mb1_FB2_BB2_IO_030,
    input wire        mb1_FB1_TB0_IO_021_mb1_FB2_BB2_IO_031,
    input wire        mb1_FB1_TB0_IO_022_mb1_FB2_BB2_IO_008,
    input wire        mb1_FB1_TB0_IO_023_mb1_FB2_BB2_IO_009,
    input wire        mb1_FB1_TB0_IO_024_mb1_FB2_BB2_IO_026,
    input wire        mb1_FB1_TB0_IO_025_mb1_FB2_BB2_IO_027,
    input wire        mb1_FB1_TB0_IO_026_mb1_FB2_BB2_IO_024,
    input wire        mb1_FB1_TB0_IO_027_mb1_FB2_BB2_IO_025,
    input wire        mb1_FB1_TB0_IO_028_mb1_FB2_BB2_IO_042,
    input wire        mb1_FB1_TB0_IO_029_mb1_FB2_BB2_IO_043,
    input wire        mb1_FB1_TB0_IO_030_mb1_FB2_BB2_IO_020,
    input wire        mb1_FB1_TB0_IO_031_mb1_FB2_BB2_IO_021,
    input wire        mb1_FB1_TB0_IO_032_mb1_FB2_BB2_IO_018,
    input wire        mb1_FB1_TB0_IO_033_mb1_FB2_BB2_IO_019,
    input wire        mb1_FB1_TB0_IO_034_mb1_FB2_BB2_IO_036,
    input wire        mb1_FB1_TB0_IO_035_mb1_FB2_BB2_IO_037,
    input wire        mb1_FB1_TB0_IO_036_mb1_FB2_BB2_IO_034,
    input wire        mb1_FB1_TB0_IO_037_mb1_FB2_BB2_IO_035,
    input wire        mb1_FB1_TB0_IO_038_mb1_FB2_BB2_IO_052,
    input wire        mb1_FB1_TB0_IO_039_mb1_FB2_BB2_IO_053,
    input wire        mb1_FB1_TB0_IO_040_mb1_FB2_BB2_IO_050,
    input wire        mb1_FB1_TB0_IO_041_mb1_FB2_BB2_IO_051,
    input wire        mb1_FB1_TB0_IO_042_mb1_FB2_BB2_IO_028,
    input wire        mb1_FB1_TB0_IO_043_mb1_FB2_BB2_IO_029,
    input wire        mb1_FB1_TB0_IO_044_mb1_FB2_BB2_IO_046,
    input wire        mb1_FB1_TB0_IO_045_mb1_FB2_BB2_IO_047,
    input wire        mb1_FB1_TB0_IO_046_mb1_FB2_BB2_IO_044,
    input wire        mb1_FB1_TB0_IO_047_mb1_FB2_BB2_IO_045,
    input wire        mb1_FB1_TB0_IO_048_mb1_FB2_BB2_IO_062,
    input wire        mb1_FB1_TB0_IO_049_mb1_FB2_BB2_IO_063,
    input wire        mb1_FB1_TB0_IO_050_mb1_FB2_BB2_IO_040,
    input wire        mb1_FB1_TB0_IO_051_mb1_FB2_BB2_IO_041,
    input wire        mb1_FB1_TB0_IO_052_mb1_FB2_BB2_IO_038,
    input wire        mb1_FB1_TB0_IO_053_mb1_FB2_BB2_IO_039,
    input wire        mb1_FB1_TB0_IO_054_mb1_FB2_BB2_IO_056,
    input wire        mb1_FB1_TB0_IO_055_mb1_FB2_BB2_IO_057,
    input wire        mb1_FB1_TB0_IO_056_mb1_FB2_BB2_IO_054,
    input wire        mb1_FB1_TB0_IO_057_mb1_FB2_BB2_IO_055,
    input wire        mb1_FB1_TB0_IO_058_mb1_FB2_BB2_IO_072,
    input wire        mb1_FB1_TB0_IO_059_mb1_FB2_BB2_IO_073,
    input wire        mb1_FB1_TB0_IO_060_mb1_FB2_BB2_IO_070,
    input wire        mb1_FB1_TB0_IO_061_mb1_FB2_BB2_IO_071,
    input wire        mb1_FB1_TB0_IO_062_mb1_FB2_BB2_IO_048,
    input wire        mb1_FB1_TB0_IO_063_mb1_FB2_BB2_IO_049,
    input wire        mb1_FB1_TB0_IO_064_mb1_FB2_BB2_IO_066,
    input wire        mb1_FB1_TB0_IO_065_mb1_FB2_BB2_IO_067,
    input wire        mb1_FB1_TB0_IO_066_mb1_FB2_BB2_IO_064,
    input wire        mb1_FB1_TB0_IO_067_mb1_FB2_BB2_IO_065,
    input wire        mb1_FB1_TB0_IO_068_mb1_FB2_BB2_IO_082,
    input wire        mb1_FB1_TB0_IO_069_mb1_FB2_BB2_IO_083,
    input wire        mb1_FB1_TB0_IO_070_mb1_FB2_BB2_IO_060,
    input wire        mb1_FB1_TB0_IO_071_mb1_FB2_BB2_IO_061,
    input wire        mb1_FB1_TB0_IO_072_mb1_FB2_BB2_IO_058,
    input wire        mb1_FB1_TB0_IO_073_mb1_FB2_BB2_IO_059,
    input wire        mb1_FB1_TB0_IO_074_mb1_FB2_BB2_IO_076,
    input wire        mb1_FB1_TB0_IO_075_mb1_FB2_BB2_IO_077,
    input wire        mb1_FB1_TB0_IO_076_mb1_FB2_BB2_IO_074,
    input wire        mb1_FB1_TB0_IO_077_mb1_FB2_BB2_IO_075,
    input wire        mb1_FB1_TB0_IO_078_mb1_FB2_BB2_IO_092,
    input wire        mb1_FB1_TB0_IO_079_mb1_FB2_BB2_IO_093,
    input wire        mb1_FB1_TB0_IO_080_mb1_FB2_BB2_IO_090,
    input wire        mb1_FB1_TB0_IO_081_mb1_FB2_BB2_IO_091,
    input wire        mb1_FB1_TB0_IO_082_mb1_FB2_BB2_IO_068,
    input wire        mb1_FB1_TB0_IO_083_mb1_FB2_BB2_IO_069,
    input wire        mb1_FB1_TB0_IO_084_mb1_FB2_BB2_IO_086,
    input wire        mb1_FB1_TB0_IO_085_mb1_FB2_BB2_IO_087,
    input wire        mb1_FB1_TB0_IO_086_mb1_FB2_BB2_IO_084,
    input wire        mb1_FB1_TB0_IO_087_mb1_FB2_BB2_IO_085,
    input wire        mb1_FB1_TB0_IO_088_mb1_FB2_BB2_IO_102,
    input wire        mb1_FB1_TB0_IO_089_mb1_FB2_BB2_IO_103,
    input wire        mb1_FB1_TB0_IO_090_mb1_FB2_BB2_IO_080,
    input wire        mb1_FB1_TB0_IO_091_mb1_FB2_BB2_IO_081,
    input wire        mb1_FB1_TB0_IO_092_mb1_FB2_BB2_IO_078,
    input wire        mb1_FB1_TB0_IO_093_mb1_FB2_BB2_IO_079,
    input wire        mb1_FB1_TB0_IO_094_mb1_FB2_BB2_IO_096,
    input wire        mb1_FB1_TB0_IO_095_mb1_FB2_BB2_IO_097,
    input wire        mb1_FB1_TB0_IO_096_mb1_FB2_BB2_IO_094,
    input wire        mb1_FB1_TB0_IO_097_mb1_FB2_BB2_IO_095,
    input wire        mb1_FB1_TB0_IO_098_mb1_FB2_BB2_IO_112,
    input wire        mb1_FB1_TB0_IO_099_mb1_FB2_BB2_IO_113,
    input wire        mb1_FB1_TB0_IO_100_mb1_FB2_BB2_IO_110,
    input wire        mb1_FB1_TB0_IO_101_mb1_FB2_BB2_IO_111,
    input wire        mb1_FB1_TB0_IO_102_mb1_FB2_BB2_IO_088,
    input wire        mb1_FB1_TB0_IO_103_mb1_FB2_BB2_IO_089,
    input wire        mb1_FB1_TB0_IO_104_mb1_FB2_BB2_IO_106,
    input wire        mb1_FB1_TB0_IO_105_mb1_FB2_BB2_IO_107,
    input wire        mb1_FB1_TB0_IO_106_mb1_FB2_BB2_IO_104,
    input wire        mb1_FB1_TB0_IO_107_mb1_FB2_BB2_IO_105,
    input wire        mb1_FB1_TB0_IO_108_mb1_FB2_BB2_IO_122,
    input wire        mb1_FB1_TB0_IO_109_mb1_FB2_BB2_IO_123,
    input wire        mb1_FB1_TB0_IO_110_mb1_FB2_BB2_IO_100,
    input wire        mb1_FB1_TB0_IO_111_mb1_FB2_BB2_IO_101,
    input wire        mb1_FB1_TB0_IO_112_mb1_FB2_BB2_IO_098,
    input wire        mb1_FB1_TB0_IO_113_mb1_FB2_BB2_IO_099,
    input wire        mb1_FB1_TB0_IO_114_mb1_FB2_BB2_IO_116,
    input wire        mb1_FB1_TB0_IO_115_mb1_FB2_BB2_IO_117,
    input wire        mb1_FB1_TB0_IO_116_mb1_FB2_BB2_IO_114,
    input wire        mb1_FB1_TB0_IO_117_mb1_FB2_BB2_IO_115,
    input wire        mb1_FB1_TB0_IO_118_mb1_FB2_BB2_IO_132,
    input wire        mb1_FB1_TB0_IO_119_mb1_FB2_BB2_IO_133,
    input wire        mb1_FB1_TB0_IO_120_mb1_FB2_BB2_IO_130,
    input wire        mb1_FB1_TB0_IO_121_mb1_FB2_BB2_IO_131,
    input wire        mb1_FB1_TB0_IO_122_mb1_FB2_BB2_IO_108,
    input wire        mb1_FB1_TB0_IO_123_mb1_FB2_BB2_IO_109,
    input wire        mb1_FB1_TB0_IO_124_mb1_FB2_BB2_IO_126,
    input wire        mb1_FB1_TB0_IO_125_mb1_FB2_BB2_IO_127,
    input wire        mb1_FB1_TB0_IO_126_mb1_FB2_BB2_IO_124,
    input wire        mb1_FB1_TB0_IO_127_mb1_FB2_BB2_IO_125,
    input wire        mb1_FB1_TB0_IO_130_mb1_FB2_BB2_IO_120,
    input wire        mb1_FB1_TB0_IO_131_mb1_FB2_BB2_IO_121,
    input wire        mb1_FB1_TB0_IO_132_mb1_FB2_BB2_IO_118,
    input wire        mb1_FB1_TB0_IO_133_mb1_FB2_BB2_IO_119,
    input wire        mb1_FB1_TB0_IO_134_mb1_FB2_BB2_IO_136,
    input wire        mb1_FB1_TB0_IO_136_mb1_FB2_BB2_IO_134);

  localparam TX_PINS            = 0;
  localparam RX_PINS            = 1460;
  localparam USE_CLK_INPUT_BUFG = 0;

  wire [RX_PINS-1:0] rx_pin;

  assign rx_pin[0] = mb1_FA2_TA0_CLKIO_N_0_mb1_FB2_TA2_CLKIO_N_7;
  assign rx_pin[1] = mb1_FA2_TA0_CLKIO_N_1_mb1_FB2_TA2_CLKIO_N_6;
  assign rx_pin[2] = mb1_FA2_TA0_CLKIO_N_2_mb1_FB2_TA2_CLKIO_N_4;
  assign rx_pin[3] = mb1_FA2_TA0_CLKIO_N_3_mb1_FB2_TA2_CLKIO_N_3;
  assign rx_pin[4] = mb1_FA2_TA0_CLKIO_N_4_mb1_FB2_TA2_CLKIO_N_2;
  assign rx_pin[5] = mb1_FA2_TA0_CLKIO_N_5_mb1_FB2_TA2_IO_010;
  assign rx_pin[6] = mb1_FA2_TA0_CLKIO_N_6_mb1_FB2_TA2_CLKIO_N_1;
  assign rx_pin[7] = mb1_FA2_TA0_CLKIO_N_7_mb1_FB2_TA2_CLKIO_N_0;
  assign rx_pin[8] = mb1_FA2_TA0_CLKIO_P_0_mb1_FB2_TA2_CLKIO_P_7;
  assign rx_pin[9] = mb1_FA2_TA0_CLKIO_P_1_mb1_FB2_TA2_CLKIO_P_6;
  assign rx_pin[10] = mb1_FA2_TA0_CLKIO_P_2_mb1_FB2_TA2_CLKIO_P_4;
  assign rx_pin[11] = mb1_FA2_TA0_CLKIO_P_3_mb1_FB2_TA2_CLKIO_P_3;
  assign rx_pin[12] = mb1_FA2_TA0_CLKIO_P_4_mb1_FB2_TA2_CLKIO_P_2;
  assign rx_pin[13] = mb1_FA2_TA0_CLKIO_P_5_mb1_FB2_TA2_IO_011;
  assign rx_pin[14] = mb1_FA2_TA0_CLKIO_P_6_mb1_FB2_TA2_CLKIO_P_1;
  assign rx_pin[15] = mb1_FA2_TA0_CLKIO_P_7_mb1_FB2_TA2_CLKIO_P_0;
  assign rx_pin[16] = mb1_FA2_TA0_IO_004_mb1_FB2_TA2_IO_006;
  assign rx_pin[17] = mb1_FA2_TA0_IO_005_mb1_FB2_TA2_IO_007;
  assign rx_pin[18] = mb1_FA2_TA0_IO_006_mb1_FB2_TA2_IO_004;
  assign rx_pin[19] = mb1_FA2_TA0_IO_007_mb1_FB2_TA2_IO_005;
  assign rx_pin[20] = mb1_FA2_TA0_IO_008_mb1_FB2_TA2_IO_022;
  assign rx_pin[21] = mb1_FA2_TA0_IO_009_mb1_FB2_TA2_IO_023;
  assign rx_pin[22] = mb1_FA2_TA0_IO_010_mb1_FB2_TA2_CLKIO_N_5;
  assign rx_pin[23] = mb1_FA2_TA0_IO_011_mb1_FB2_TA2_CLKIO_P_5;
  assign rx_pin[24] = mb1_FA2_TA0_IO_012_mb1_FB2_TA2_IO_012;
  assign rx_pin[25] = mb1_FA2_TA0_IO_013_mb1_FB2_TA2_IO_013;
  assign rx_pin[26] = mb1_FA2_TA0_IO_014_mb1_FB2_TA2_IO_016;
  assign rx_pin[27] = mb1_FA2_TA0_IO_015_mb1_FB2_TA2_IO_017;
  assign rx_pin[28] = mb1_FA2_TA0_IO_016_mb1_FB2_TA2_IO_014;
  assign rx_pin[29] = mb1_FA2_TA0_IO_017_mb1_FB2_TA2_IO_015;
  assign rx_pin[30] = mb1_FA2_TA0_IO_018_mb1_FB2_TA2_IO_032;
  assign rx_pin[31] = mb1_FA2_TA0_IO_019_mb1_FB2_TA2_IO_033;
  assign rx_pin[32] = mb1_FA2_TA0_IO_020_mb1_FB2_TA2_IO_030;
  assign rx_pin[33] = mb1_FA2_TA0_IO_021_mb1_FB2_TA2_IO_031;
  assign rx_pin[34] = mb1_FA2_TA0_IO_022_mb1_FB2_TA2_IO_008;
  assign rx_pin[35] = mb1_FA2_TA0_IO_023_mb1_FB2_TA2_IO_009;
  assign rx_pin[36] = mb1_FA2_TA0_IO_024_mb1_FB2_TA2_IO_026;
  assign rx_pin[37] = mb1_FA2_TA0_IO_025_mb1_FB2_TA2_IO_027;
  assign rx_pin[38] = mb1_FA2_TA0_IO_026_mb1_FB2_TA2_IO_024;
  assign rx_pin[39] = mb1_FA2_TA0_IO_027_mb1_FB2_TA2_IO_025;
  assign rx_pin[40] = mb1_FA2_TA0_IO_028_mb1_FB2_TA2_IO_042;
  assign rx_pin[41] = mb1_FA2_TA0_IO_029_mb1_FB2_TA2_IO_043;
  assign rx_pin[42] = mb1_FA2_TA0_IO_030_mb1_FB2_TA2_IO_020;
  assign rx_pin[43] = mb1_FA2_TA0_IO_031_mb1_FB2_TA2_IO_021;
  assign rx_pin[44] = mb1_FA2_TA0_IO_032_mb1_FB2_TA2_IO_018;
  assign rx_pin[45] = mb1_FA2_TA0_IO_033_mb1_FB2_TA2_IO_019;
  assign rx_pin[46] = mb1_FA2_TA0_IO_034_mb1_FB2_TA2_IO_036;
  assign rx_pin[47] = mb1_FA2_TA0_IO_035_mb1_FB2_TA2_IO_037;
  assign rx_pin[48] = mb1_FA2_TA0_IO_036_mb1_FB2_TA2_IO_034;
  assign rx_pin[49] = mb1_FA2_TA0_IO_037_mb1_FB2_TA2_IO_035;
  assign rx_pin[50] = mb1_FA2_TA0_IO_038_mb1_FB2_TA2_IO_052;
  assign rx_pin[51] = mb1_FA2_TA0_IO_039_mb1_FB2_TA2_IO_053;
  assign rx_pin[52] = mb1_FA2_TA0_IO_040_mb1_FB2_TA2_IO_050;
  assign rx_pin[53] = mb1_FA2_TA0_IO_041_mb1_FB2_TA2_IO_051;
  assign rx_pin[54] = mb1_FA2_TA0_IO_042_mb1_FB2_TA2_IO_028;
  assign rx_pin[55] = mb1_FA2_TA0_IO_043_mb1_FB2_TA2_IO_029;
  assign rx_pin[56] = mb1_FA2_TA0_IO_044_mb1_FB2_TA2_IO_046;
  assign rx_pin[57] = mb1_FA2_TA0_IO_045_mb1_FB2_TA2_IO_047;
  assign rx_pin[58] = mb1_FA2_TA0_IO_046_mb1_FB2_TA2_IO_044;
  assign rx_pin[59] = mb1_FA2_TA0_IO_047_mb1_FB2_TA2_IO_045;
  assign rx_pin[60] = mb1_FA2_TA0_IO_048_mb1_FB2_TA2_IO_062;
  assign rx_pin[61] = mb1_FA2_TA0_IO_049_mb1_FB2_TA2_IO_063;
  assign rx_pin[62] = mb1_FA2_TA0_IO_050_mb1_FB2_TA2_IO_040;
  assign rx_pin[63] = mb1_FA2_TA0_IO_051_mb1_FB2_TA2_IO_041;
  assign rx_pin[64] = mb1_FA2_TA0_IO_052_mb1_FB2_TA2_IO_038;
  assign rx_pin[65] = mb1_FA2_TA0_IO_053_mb1_FB2_TA2_IO_039;
  assign rx_pin[66] = mb1_FA2_TA0_IO_054_mb1_FB2_TA2_IO_056;
  assign rx_pin[67] = mb1_FA2_TA0_IO_055_mb1_FB2_TA2_IO_057;
  assign rx_pin[68] = mb1_FA2_TA0_IO_056_mb1_FB2_TA2_IO_054;
  assign rx_pin[69] = mb1_FA2_TA0_IO_057_mb1_FB2_TA2_IO_055;
  assign rx_pin[70] = mb1_FA2_TA0_IO_058_mb1_FB2_TA2_IO_072;
  assign rx_pin[71] = mb1_FA2_TA0_IO_059_mb1_FB2_TA2_IO_073;
  assign rx_pin[72] = mb1_FA2_TA0_IO_060_mb1_FB2_TA2_IO_070;
  assign rx_pin[73] = mb1_FA2_TA0_IO_061_mb1_FB2_TA2_IO_071;
  assign rx_pin[74] = mb1_FA2_TA0_IO_062_mb1_FB2_TA2_IO_048;
  assign rx_pin[75] = mb1_FA2_TA0_IO_063_mb1_FB2_TA2_IO_049;
  assign rx_pin[76] = mb1_FA2_TA0_IO_064_mb1_FB2_TA2_IO_066;
  assign rx_pin[77] = mb1_FA2_TA0_IO_065_mb1_FB2_TA2_IO_067;
  assign rx_pin[78] = mb1_FA2_TA0_IO_066_mb1_FB2_TA2_IO_064;
  assign rx_pin[79] = mb1_FA2_TA0_IO_067_mb1_FB2_TA2_IO_065;
  assign rx_pin[80] = mb1_FA2_TA0_IO_068_mb1_FB2_TA2_IO_082;
  assign rx_pin[81] = mb1_FA2_TA0_IO_069_mb1_FB2_TA2_IO_083;
  assign rx_pin[82] = mb1_FA2_TA0_IO_070_mb1_FB2_TA2_IO_060;
  assign rx_pin[83] = mb1_FA2_TA0_IO_071_mb1_FB2_TA2_IO_061;
  assign rx_pin[84] = mb1_FA2_TA0_IO_072_mb1_FB2_TA2_IO_058;
  assign rx_pin[85] = mb1_FA2_TA0_IO_073_mb1_FB2_TA2_IO_059;
  assign rx_pin[86] = mb1_FA2_TA0_IO_074_mb1_FB2_TA2_IO_076;
  assign rx_pin[87] = mb1_FA2_TA0_IO_075_mb1_FB2_TA2_IO_077;
  assign rx_pin[88] = mb1_FA2_TA0_IO_076_mb1_FB2_TA2_IO_074;
  assign rx_pin[89] = mb1_FA2_TA0_IO_077_mb1_FB2_TA2_IO_075;
  assign rx_pin[90] = mb1_FA2_TA0_IO_078_mb1_FB2_TA2_IO_092;
  assign rx_pin[91] = mb1_FA2_TA0_IO_079_mb1_FB2_TA2_IO_093;
  assign rx_pin[92] = mb1_FA2_TA0_IO_080_mb1_FB2_TA2_IO_090;
  assign rx_pin[93] = mb1_FA2_TA0_IO_081_mb1_FB2_TA2_IO_091;
  assign rx_pin[94] = mb1_FA2_TA0_IO_082_mb1_FB2_TA2_IO_068;
  assign rx_pin[95] = mb1_FA2_TA0_IO_083_mb1_FB2_TA2_IO_069;
  assign rx_pin[96] = mb1_FA2_TA0_IO_084_mb1_FB2_TA2_IO_086;
  assign rx_pin[97] = mb1_FA2_TA0_IO_085_mb1_FB2_TA2_IO_087;
  assign rx_pin[98] = mb1_FA2_TA0_IO_086_mb1_FB2_TA2_IO_084;
  assign rx_pin[99] = mb1_FA2_TA0_IO_087_mb1_FB2_TA2_IO_085;
  assign rx_pin[100] = mb1_FA2_TA0_IO_088_mb1_FB2_TA2_IO_102;
  assign rx_pin[101] = mb1_FA2_TA0_IO_089_mb1_FB2_TA2_IO_103;
  assign rx_pin[102] = mb1_FA2_TA0_IO_090_mb1_FB2_TA2_IO_080;
  assign rx_pin[103] = mb1_FA2_TA0_IO_091_mb1_FB2_TA2_IO_081;
  assign rx_pin[104] = mb1_FA2_TA0_IO_092_mb1_FB2_TA2_IO_078;
  assign rx_pin[105] = mb1_FA2_TA0_IO_093_mb1_FB2_TA2_IO_079;
  assign rx_pin[106] = mb1_FA2_TA0_IO_094_mb1_FB2_TA2_IO_096;
  assign rx_pin[107] = mb1_FA2_TA0_IO_095_mb1_FB2_TA2_IO_097;
  assign rx_pin[108] = mb1_FA2_TA0_IO_096_mb1_FB2_TA2_IO_094;
  assign rx_pin[109] = mb1_FA2_TA0_IO_097_mb1_FB2_TA2_IO_095;
  assign rx_pin[110] = mb1_FA2_TA0_IO_098_mb1_FB2_TA2_IO_112;
  assign rx_pin[111] = mb1_FA2_TA0_IO_099_mb1_FB2_TA2_IO_113;
  assign rx_pin[112] = mb1_FA2_TA0_IO_100_mb1_FB2_TA2_IO_110;
  assign rx_pin[113] = mb1_FA2_TA0_IO_101_mb1_FB2_TA2_IO_111;
  assign rx_pin[114] = mb1_FA2_TA0_IO_102_mb1_FB2_TA2_IO_088;
  assign rx_pin[115] = mb1_FA2_TA0_IO_103_mb1_FB2_TA2_IO_089;
  assign rx_pin[116] = mb1_FA2_TA0_IO_104_mb1_FB2_TA2_IO_106;
  assign rx_pin[117] = mb1_FA2_TA0_IO_105_mb1_FB2_TA2_IO_107;
  assign rx_pin[118] = mb1_FA2_TA0_IO_106_mb1_FB2_TA2_IO_104;
  assign rx_pin[119] = mb1_FA2_TA0_IO_107_mb1_FB2_TA2_IO_105;
  assign rx_pin[120] = mb1_FA2_TA0_IO_108_mb1_FB2_TA2_IO_122;
  assign rx_pin[121] = mb1_FA2_TA0_IO_109_mb1_FB2_TA2_IO_123;
  assign rx_pin[122] = mb1_FA2_TA0_IO_110_mb1_FB2_TA2_IO_100;
  assign rx_pin[123] = mb1_FA2_TA0_IO_111_mb1_FB2_TA2_IO_101;
  assign rx_pin[124] = mb1_FA2_TA0_IO_112_mb1_FB2_TA2_IO_098;
  assign rx_pin[125] = mb1_FA2_TA0_IO_113_mb1_FB2_TA2_IO_099;
  assign rx_pin[126] = mb1_FA2_TA0_IO_114_mb1_FB2_TA2_IO_116;
  assign rx_pin[127] = mb1_FA2_TA0_IO_115_mb1_FB2_TA2_IO_117;
  assign rx_pin[128] = mb1_FA2_TA0_IO_116_mb1_FB2_TA2_IO_114;
  assign rx_pin[129] = mb1_FA2_TA0_IO_117_mb1_FB2_TA2_IO_115;
  assign rx_pin[130] = mb1_FA2_TA0_IO_118_mb1_FB2_TA2_IO_132;
  assign rx_pin[131] = mb1_FA2_TA0_IO_119_mb1_FB2_TA2_IO_133;
  assign rx_pin[132] = mb1_FA2_TA0_IO_120_mb1_FB2_TA2_IO_130;
  assign rx_pin[133] = mb1_FA2_TA0_IO_121_mb1_FB2_TA2_IO_131;
  assign rx_pin[134] = mb1_FA2_TA0_IO_122_mb1_FB2_TA2_IO_108;
  assign rx_pin[135] = mb1_FA2_TA0_IO_123_mb1_FB2_TA2_IO_109;
  assign rx_pin[136] = mb1_FA2_TA0_IO_124_mb1_FB2_TA2_IO_126;
  assign rx_pin[137] = mb1_FA2_TA0_IO_125_mb1_FB2_TA2_IO_127;
  assign rx_pin[138] = mb1_FA2_TA0_IO_126_mb1_FB2_TA2_IO_124;
  assign rx_pin[139] = mb1_FA2_TA0_IO_127_mb1_FB2_TA2_IO_125;
  assign rx_pin[140] = mb1_FA2_TA0_IO_130_mb1_FB2_TA2_IO_120;
  assign rx_pin[141] = mb1_FA2_TA0_IO_131_mb1_FB2_TA2_IO_121;
  assign rx_pin[142] = mb1_FA2_TA0_IO_132_mb1_FB2_TA2_IO_118;
  assign rx_pin[143] = mb1_FA2_TA0_IO_133_mb1_FB2_TA2_IO_119;
  assign rx_pin[144] = mb1_FA2_TA0_IO_134_mb1_FB2_TA2_IO_136;
  assign rx_pin[145] = mb1_FA2_TA0_IO_136_mb1_FB2_TA2_IO_134;
  assign rx_pin[146] = mb1_FA2_BA0_CLKIO_N_0_mb1_FB2_TB0_CLKIO_N_7;
  assign rx_pin[147] = mb1_FA2_BA0_CLKIO_N_1_mb1_FB2_TB0_CLKIO_N_6;
  assign rx_pin[148] = mb1_FA2_BA0_CLKIO_N_2_mb1_FB2_TB0_CLKIO_N_4;
  assign rx_pin[149] = mb1_FA2_BA0_CLKIO_N_3_mb1_FB2_TB0_CLKIO_N_3;
  assign rx_pin[150] = mb1_FA2_BA0_CLKIO_N_4_mb1_FB2_TB0_CLKIO_N_2;
  assign rx_pin[151] = mb1_FA2_BA0_CLKIO_N_5_mb1_FB2_TB0_IO_010;
  assign rx_pin[152] = mb1_FA2_BA0_CLKIO_N_6_mb1_FB2_TB0_CLKIO_N_1;
  assign rx_pin[153] = mb1_FA2_BA0_CLKIO_N_7_mb1_FB2_TB0_CLKIO_N_0;
  assign rx_pin[154] = mb1_FA2_BA0_CLKIO_P_0_mb1_FB2_TB0_CLKIO_P_7;
  assign rx_pin[155] = mb1_FA2_BA0_CLKIO_P_1_mb1_FB2_TB0_CLKIO_P_6;
  assign rx_pin[156] = mb1_FA2_BA0_CLKIO_P_2_mb1_FB2_TB0_CLKIO_P_4;
  assign rx_pin[157] = mb1_FA2_BA0_CLKIO_P_3_mb1_FB2_TB0_CLKIO_P_3;
  assign rx_pin[158] = mb1_FA2_BA0_CLKIO_P_4_mb1_FB2_TB0_CLKIO_P_2;
  assign rx_pin[159] = mb1_FA2_BA0_CLKIO_P_5_mb1_FB2_TB0_IO_011;
  assign rx_pin[160] = mb1_FA2_BA0_CLKIO_P_6_mb1_FB2_TB0_CLKIO_P_1;
  assign rx_pin[161] = mb1_FA2_BA0_CLKIO_P_7_mb1_FB2_TB0_CLKIO_P_0;
  assign rx_pin[162] = mb1_FA2_BA0_IO_004_mb1_FB2_TB0_IO_006;
  assign rx_pin[163] = mb1_FA2_BA0_IO_005_mb1_FB2_TB0_IO_007;
  assign rx_pin[164] = mb1_FA2_BA0_IO_006_mb1_FB2_TB0_IO_004;
  assign rx_pin[165] = mb1_FA2_BA0_IO_007_mb1_FB2_TB0_IO_005;
  assign rx_pin[166] = mb1_FA2_BA0_IO_008_mb1_FB2_TB0_IO_022;
  assign rx_pin[167] = mb1_FA2_BA0_IO_009_mb1_FB2_TB0_IO_023;
  assign rx_pin[168] = mb1_FA2_BA0_IO_010_mb1_FB2_TB0_CLKIO_N_5;
  assign rx_pin[169] = mb1_FA2_BA0_IO_011_mb1_FB2_TB0_CLKIO_P_5;
  assign rx_pin[170] = mb1_FA2_BA0_IO_012_mb1_FB2_TB0_IO_012;
  assign rx_pin[171] = mb1_FA2_BA0_IO_013_mb1_FB2_TB0_IO_013;
  assign rx_pin[172] = mb1_FA2_BA0_IO_014_mb1_FB2_TB0_IO_016;
  assign rx_pin[173] = mb1_FA2_BA0_IO_015_mb1_FB2_TB0_IO_017;
  assign rx_pin[174] = mb1_FA2_BA0_IO_016_mb1_FB2_TB0_IO_014;
  assign rx_pin[175] = mb1_FA2_BA0_IO_017_mb1_FB2_TB0_IO_015;
  assign rx_pin[176] = mb1_FA2_BA0_IO_018_mb1_FB2_TB0_IO_032;
  assign rx_pin[177] = mb1_FA2_BA0_IO_019_mb1_FB2_TB0_IO_033;
  assign rx_pin[178] = mb1_FA2_BA0_IO_020_mb1_FB2_TB0_IO_030;
  assign rx_pin[179] = mb1_FA2_BA0_IO_021_mb1_FB2_TB0_IO_031;
  assign rx_pin[180] = mb1_FA2_BA0_IO_022_mb1_FB2_TB0_IO_008;
  assign rx_pin[181] = mb1_FA2_BA0_IO_023_mb1_FB2_TB0_IO_009;
  assign rx_pin[182] = mb1_FA2_BA0_IO_024_mb1_FB2_TB0_IO_026;
  assign rx_pin[183] = mb1_FA2_BA0_IO_025_mb1_FB2_TB0_IO_027;
  assign rx_pin[184] = mb1_FA2_BA0_IO_026_mb1_FB2_TB0_IO_024;
  assign rx_pin[185] = mb1_FA2_BA0_IO_027_mb1_FB2_TB0_IO_025;
  assign rx_pin[186] = mb1_FA2_BA0_IO_028_mb1_FB2_TB0_IO_042;
  assign rx_pin[187] = mb1_FA2_BA0_IO_029_mb1_FB2_TB0_IO_043;
  assign rx_pin[188] = mb1_FA2_BA0_IO_030_mb1_FB2_TB0_IO_020;
  assign rx_pin[189] = mb1_FA2_BA0_IO_031_mb1_FB2_TB0_IO_021;
  assign rx_pin[190] = mb1_FA2_BA0_IO_032_mb1_FB2_TB0_IO_018;
  assign rx_pin[191] = mb1_FA2_BA0_IO_033_mb1_FB2_TB0_IO_019;
  assign rx_pin[192] = mb1_FA2_BA0_IO_034_mb1_FB2_TB0_IO_036;
  assign rx_pin[193] = mb1_FA2_BA0_IO_035_mb1_FB2_TB0_IO_037;
  assign rx_pin[194] = mb1_FA2_BA0_IO_036_mb1_FB2_TB0_IO_034;
  assign rx_pin[195] = mb1_FA2_BA0_IO_037_mb1_FB2_TB0_IO_035;
  assign rx_pin[196] = mb1_FA2_BA0_IO_038_mb1_FB2_TB0_IO_052;
  assign rx_pin[197] = mb1_FA2_BA0_IO_039_mb1_FB2_TB0_IO_053;
  assign rx_pin[198] = mb1_FA2_BA0_IO_040_mb1_FB2_TB0_IO_050;
  assign rx_pin[199] = mb1_FA2_BA0_IO_041_mb1_FB2_TB0_IO_051;
  assign rx_pin[200] = mb1_FA2_BA0_IO_042_mb1_FB2_TB0_IO_028;
  assign rx_pin[201] = mb1_FA2_BA0_IO_043_mb1_FB2_TB0_IO_029;
  assign rx_pin[202] = mb1_FA2_BA0_IO_044_mb1_FB2_TB0_IO_046;
  assign rx_pin[203] = mb1_FA2_BA0_IO_045_mb1_FB2_TB0_IO_047;
  assign rx_pin[204] = mb1_FA2_BA0_IO_046_mb1_FB2_TB0_IO_044;
  assign rx_pin[205] = mb1_FA2_BA0_IO_047_mb1_FB2_TB0_IO_045;
  assign rx_pin[206] = mb1_FA2_BA0_IO_048_mb1_FB2_TB0_IO_062;
  assign rx_pin[207] = mb1_FA2_BA0_IO_049_mb1_FB2_TB0_IO_063;
  assign rx_pin[208] = mb1_FA2_BA0_IO_050_mb1_FB2_TB0_IO_040;
  assign rx_pin[209] = mb1_FA2_BA0_IO_051_mb1_FB2_TB0_IO_041;
  assign rx_pin[210] = mb1_FA2_BA0_IO_052_mb1_FB2_TB0_IO_038;
  assign rx_pin[211] = mb1_FA2_BA0_IO_053_mb1_FB2_TB0_IO_039;
  assign rx_pin[212] = mb1_FA2_BA0_IO_054_mb1_FB2_TB0_IO_056;
  assign rx_pin[213] = mb1_FA2_BA0_IO_055_mb1_FB2_TB0_IO_057;
  assign rx_pin[214] = mb1_FA2_BA0_IO_056_mb1_FB2_TB0_IO_054;
  assign rx_pin[215] = mb1_FA2_BA0_IO_057_mb1_FB2_TB0_IO_055;
  assign rx_pin[216] = mb1_FA2_BA0_IO_058_mb1_FB2_TB0_IO_072;
  assign rx_pin[217] = mb1_FA2_BA0_IO_059_mb1_FB2_TB0_IO_073;
  assign rx_pin[218] = mb1_FA2_BA0_IO_060_mb1_FB2_TB0_IO_070;
  assign rx_pin[219] = mb1_FA2_BA0_IO_061_mb1_FB2_TB0_IO_071;
  assign rx_pin[220] = mb1_FA2_BA0_IO_062_mb1_FB2_TB0_IO_048;
  assign rx_pin[221] = mb1_FA2_BA0_IO_063_mb1_FB2_TB0_IO_049;
  assign rx_pin[222] = mb1_FA2_BA0_IO_064_mb1_FB2_TB0_IO_066;
  assign rx_pin[223] = mb1_FA2_BA0_IO_065_mb1_FB2_TB0_IO_067;
  assign rx_pin[224] = mb1_FA2_BA0_IO_066_mb1_FB2_TB0_IO_064;
  assign rx_pin[225] = mb1_FA2_BA0_IO_067_mb1_FB2_TB0_IO_065;
  assign rx_pin[226] = mb1_FA2_BA0_IO_068_mb1_FB2_TB0_IO_082;
  assign rx_pin[227] = mb1_FA2_BA0_IO_069_mb1_FB2_TB0_IO_083;
  assign rx_pin[228] = mb1_FA2_BA0_IO_070_mb1_FB2_TB0_IO_060;
  assign rx_pin[229] = mb1_FA2_BA0_IO_071_mb1_FB2_TB0_IO_061;
  assign rx_pin[230] = mb1_FA2_BA0_IO_072_mb1_FB2_TB0_IO_058;
  assign rx_pin[231] = mb1_FA2_BA0_IO_073_mb1_FB2_TB0_IO_059;
  assign rx_pin[232] = mb1_FA2_BA0_IO_074_mb1_FB2_TB0_IO_076;
  assign rx_pin[233] = mb1_FA2_BA0_IO_075_mb1_FB2_TB0_IO_077;
  assign rx_pin[234] = mb1_FA2_BA0_IO_076_mb1_FB2_TB0_IO_074;
  assign rx_pin[235] = mb1_FA2_BA0_IO_077_mb1_FB2_TB0_IO_075;
  assign rx_pin[236] = mb1_FA2_BA0_IO_078_mb1_FB2_TB0_IO_092;
  assign rx_pin[237] = mb1_FA2_BA0_IO_079_mb1_FB2_TB0_IO_093;
  assign rx_pin[238] = mb1_FA2_BA0_IO_080_mb1_FB2_TB0_IO_090;
  assign rx_pin[239] = mb1_FA2_BA0_IO_081_mb1_FB2_TB0_IO_091;
  assign rx_pin[240] = mb1_FA2_BA0_IO_082_mb1_FB2_TB0_IO_068;
  assign rx_pin[241] = mb1_FA2_BA0_IO_083_mb1_FB2_TB0_IO_069;
  assign rx_pin[242] = mb1_FA2_BA0_IO_084_mb1_FB2_TB0_IO_086;
  assign rx_pin[243] = mb1_FA2_BA0_IO_085_mb1_FB2_TB0_IO_087;
  assign rx_pin[244] = mb1_FA2_BA0_IO_086_mb1_FB2_TB0_IO_084;
  assign rx_pin[245] = mb1_FA2_BA0_IO_087_mb1_FB2_TB0_IO_085;
  assign rx_pin[246] = mb1_FA2_BA0_IO_088_mb1_FB2_TB0_IO_102;
  assign rx_pin[247] = mb1_FA2_BA0_IO_089_mb1_FB2_TB0_IO_103;
  assign rx_pin[248] = mb1_FA2_BA0_IO_090_mb1_FB2_TB0_IO_080;
  assign rx_pin[249] = mb1_FA2_BA0_IO_091_mb1_FB2_TB0_IO_081;
  assign rx_pin[250] = mb1_FA2_BA0_IO_092_mb1_FB2_TB0_IO_078;
  assign rx_pin[251] = mb1_FA2_BA0_IO_093_mb1_FB2_TB0_IO_079;
  assign rx_pin[252] = mb1_FA2_BA0_IO_094_mb1_FB2_TB0_IO_096;
  assign rx_pin[253] = mb1_FA2_BA0_IO_095_mb1_FB2_TB0_IO_097;
  assign rx_pin[254] = mb1_FA2_BA0_IO_096_mb1_FB2_TB0_IO_094;
  assign rx_pin[255] = mb1_FA2_BA0_IO_097_mb1_FB2_TB0_IO_095;
  assign rx_pin[256] = mb1_FA2_BA0_IO_098_mb1_FB2_TB0_IO_112;
  assign rx_pin[257] = mb1_FA2_BA0_IO_099_mb1_FB2_TB0_IO_113;
  assign rx_pin[258] = mb1_FA2_BA0_IO_100_mb1_FB2_TB0_IO_110;
  assign rx_pin[259] = mb1_FA2_BA0_IO_101_mb1_FB2_TB0_IO_111;
  assign rx_pin[260] = mb1_FA2_BA0_IO_102_mb1_FB2_TB0_IO_088;
  assign rx_pin[261] = mb1_FA2_BA0_IO_103_mb1_FB2_TB0_IO_089;
  assign rx_pin[262] = mb1_FA2_BA0_IO_104_mb1_FB2_TB0_IO_106;
  assign rx_pin[263] = mb1_FA2_BA0_IO_105_mb1_FB2_TB0_IO_107;
  assign rx_pin[264] = mb1_FA2_BA0_IO_106_mb1_FB2_TB0_IO_104;
  assign rx_pin[265] = mb1_FA2_BA0_IO_107_mb1_FB2_TB0_IO_105;
  assign rx_pin[266] = mb1_FA2_BA0_IO_108_mb1_FB2_TB0_IO_122;
  assign rx_pin[267] = mb1_FA2_BA0_IO_109_mb1_FB2_TB0_IO_123;
  assign rx_pin[268] = mb1_FA2_BA0_IO_110_mb1_FB2_TB0_IO_100;
  assign rx_pin[269] = mb1_FA2_BA0_IO_111_mb1_FB2_TB0_IO_101;
  assign rx_pin[270] = mb1_FA2_BA0_IO_112_mb1_FB2_TB0_IO_098;
  assign rx_pin[271] = mb1_FA2_BA0_IO_113_mb1_FB2_TB0_IO_099;
  assign rx_pin[272] = mb1_FA2_BA0_IO_114_mb1_FB2_TB0_IO_116;
  assign rx_pin[273] = mb1_FA2_BA0_IO_115_mb1_FB2_TB0_IO_117;
  assign rx_pin[274] = mb1_FA2_BA0_IO_116_mb1_FB2_TB0_IO_114;
  assign rx_pin[275] = mb1_FA2_BA0_IO_117_mb1_FB2_TB0_IO_115;
  assign rx_pin[276] = mb1_FA2_BA0_IO_118_mb1_FB2_TB0_IO_132;
  assign rx_pin[277] = mb1_FA2_BA0_IO_119_mb1_FB2_TB0_IO_133;
  assign rx_pin[278] = mb1_FA2_BA0_IO_120_mb1_FB2_TB0_IO_130;
  assign rx_pin[279] = mb1_FA2_BA0_IO_121_mb1_FB2_TB0_IO_131;
  assign rx_pin[280] = mb1_FA2_BA0_IO_122_mb1_FB2_TB0_IO_108;
  assign rx_pin[281] = mb1_FA2_BA0_IO_123_mb1_FB2_TB0_IO_109;
  assign rx_pin[282] = mb1_FA2_BA0_IO_124_mb1_FB2_TB0_IO_126;
  assign rx_pin[283] = mb1_FA2_BA0_IO_125_mb1_FB2_TB0_IO_127;
  assign rx_pin[284] = mb1_FA2_BA0_IO_126_mb1_FB2_TB0_IO_124;
  assign rx_pin[285] = mb1_FA2_BA0_IO_127_mb1_FB2_TB0_IO_125;
  assign rx_pin[286] = mb1_FA2_BA0_IO_130_mb1_FB2_TB0_IO_120;
  assign rx_pin[287] = mb1_FA2_BA0_IO_131_mb1_FB2_TB0_IO_121;
  assign rx_pin[288] = mb1_FA2_BA0_IO_132_mb1_FB2_TB0_IO_118;
  assign rx_pin[289] = mb1_FA2_BA0_IO_133_mb1_FB2_TB0_IO_119;
  assign rx_pin[290] = mb1_FA2_BA0_IO_134_mb1_FB2_TB0_IO_136;
  assign rx_pin[291] = mb1_FA2_BA0_IO_136_mb1_FB2_TB0_IO_134;
  assign rx_pin[292] = mb1_FA2_TA2_CLKIO_N_0_mb1_FB2_TB1_CLKIO_N_7;
  assign rx_pin[293] = mb1_FA2_TA2_CLKIO_N_1_mb1_FB2_TB1_CLKIO_N_6;
  assign rx_pin[294] = mb1_FA2_TA2_CLKIO_N_2_mb1_FB2_TB1_CLKIO_N_4;
  assign rx_pin[295] = mb1_FA2_TA2_CLKIO_N_3_mb1_FB2_TB1_CLKIO_N_3;
  assign rx_pin[296] = mb1_FA2_TA2_CLKIO_N_4_mb1_FB2_TB1_CLKIO_N_2;
  assign rx_pin[297] = mb1_FA2_TA2_CLKIO_N_5_mb1_FB2_TB1_IO_010;
  assign rx_pin[298] = mb1_FA2_TA2_CLKIO_N_6_mb1_FB2_TB1_CLKIO_N_1;
  assign rx_pin[299] = mb1_FA2_TA2_CLKIO_N_7_mb1_FB2_TB1_CLKIO_N_0;
  assign rx_pin[300] = mb1_FA2_TA2_CLKIO_P_0_mb1_FB2_TB1_CLKIO_P_7;
  assign rx_pin[301] = mb1_FA2_TA2_CLKIO_P_1_mb1_FB2_TB1_CLKIO_P_6;
  assign rx_pin[302] = mb1_FA2_TA2_CLKIO_P_2_mb1_FB2_TB1_CLKIO_P_4;
  assign rx_pin[303] = mb1_FA2_TA2_CLKIO_P_3_mb1_FB2_TB1_CLKIO_P_3;
  assign rx_pin[304] = mb1_FA2_TA2_CLKIO_P_4_mb1_FB2_TB1_CLKIO_P_2;
  assign rx_pin[305] = mb1_FA2_TA2_CLKIO_P_5_mb1_FB2_TB1_IO_011;
  assign rx_pin[306] = mb1_FA2_TA2_CLKIO_P_6_mb1_FB2_TB1_CLKIO_P_1;
  assign rx_pin[307] = mb1_FA2_TA2_CLKIO_P_7_mb1_FB2_TB1_CLKIO_P_0;
  assign rx_pin[308] = mb1_FA2_TA2_IO_004_mb1_FB2_TB1_IO_006;
  assign rx_pin[309] = mb1_FA2_TA2_IO_005_mb1_FB2_TB1_IO_007;
  assign rx_pin[310] = mb1_FA2_TA2_IO_006_mb1_FB2_TB1_IO_004;
  assign rx_pin[311] = mb1_FA2_TA2_IO_007_mb1_FB2_TB1_IO_005;
  assign rx_pin[312] = mb1_FA2_TA2_IO_008_mb1_FB2_TB1_IO_022;
  assign rx_pin[313] = mb1_FA2_TA2_IO_009_mb1_FB2_TB1_IO_023;
  assign rx_pin[314] = mb1_FA2_TA2_IO_010_mb1_FB2_TB1_CLKIO_N_5;
  assign rx_pin[315] = mb1_FA2_TA2_IO_011_mb1_FB2_TB1_CLKIO_P_5;
  assign rx_pin[316] = mb1_FA2_TA2_IO_012_mb1_FB2_TB1_IO_012;
  assign rx_pin[317] = mb1_FA2_TA2_IO_013_mb1_FB2_TB1_IO_013;
  assign rx_pin[318] = mb1_FA2_TA2_IO_014_mb1_FB2_TB1_IO_016;
  assign rx_pin[319] = mb1_FA2_TA2_IO_015_mb1_FB2_TB1_IO_017;
  assign rx_pin[320] = mb1_FA2_TA2_IO_016_mb1_FB2_TB1_IO_014;
  assign rx_pin[321] = mb1_FA2_TA2_IO_017_mb1_FB2_TB1_IO_015;
  assign rx_pin[322] = mb1_FA2_TA2_IO_018_mb1_FB2_TB1_IO_032;
  assign rx_pin[323] = mb1_FA2_TA2_IO_019_mb1_FB2_TB1_IO_033;
  assign rx_pin[324] = mb1_FA2_TA2_IO_020_mb1_FB2_TB1_IO_030;
  assign rx_pin[325] = mb1_FA2_TA2_IO_021_mb1_FB2_TB1_IO_031;
  assign rx_pin[326] = mb1_FA2_TA2_IO_022_mb1_FB2_TB1_IO_008;
  assign rx_pin[327] = mb1_FA2_TA2_IO_023_mb1_FB2_TB1_IO_009;
  assign rx_pin[328] = mb1_FA2_TA2_IO_024_mb1_FB2_TB1_IO_026;
  assign rx_pin[329] = mb1_FA2_TA2_IO_025_mb1_FB2_TB1_IO_027;
  assign rx_pin[330] = mb1_FA2_TA2_IO_026_mb1_FB2_TB1_IO_024;
  assign rx_pin[331] = mb1_FA2_TA2_IO_027_mb1_FB2_TB1_IO_025;
  assign rx_pin[332] = mb1_FA2_TA2_IO_028_mb1_FB2_TB1_IO_042;
  assign rx_pin[333] = mb1_FA2_TA2_IO_029_mb1_FB2_TB1_IO_043;
  assign rx_pin[334] = mb1_FA2_TA2_IO_030_mb1_FB2_TB1_IO_020;
  assign rx_pin[335] = mb1_FA2_TA2_IO_031_mb1_FB2_TB1_IO_021;
  assign rx_pin[336] = mb1_FA2_TA2_IO_032_mb1_FB2_TB1_IO_018;
  assign rx_pin[337] = mb1_FA2_TA2_IO_033_mb1_FB2_TB1_IO_019;
  assign rx_pin[338] = mb1_FA2_TA2_IO_034_mb1_FB2_TB1_IO_036;
  assign rx_pin[339] = mb1_FA2_TA2_IO_035_mb1_FB2_TB1_IO_037;
  assign rx_pin[340] = mb1_FA2_TA2_IO_036_mb1_FB2_TB1_IO_034;
  assign rx_pin[341] = mb1_FA2_TA2_IO_037_mb1_FB2_TB1_IO_035;
  assign rx_pin[342] = mb1_FA2_TA2_IO_038_mb1_FB2_TB1_IO_052;
  assign rx_pin[343] = mb1_FA2_TA2_IO_039_mb1_FB2_TB1_IO_053;
  assign rx_pin[344] = mb1_FA2_TA2_IO_040_mb1_FB2_TB1_IO_050;
  assign rx_pin[345] = mb1_FA2_TA2_IO_041_mb1_FB2_TB1_IO_051;
  assign rx_pin[346] = mb1_FA2_TA2_IO_042_mb1_FB2_TB1_IO_028;
  assign rx_pin[347] = mb1_FA2_TA2_IO_043_mb1_FB2_TB1_IO_029;
  assign rx_pin[348] = mb1_FA2_TA2_IO_044_mb1_FB2_TB1_IO_046;
  assign rx_pin[349] = mb1_FA2_TA2_IO_045_mb1_FB2_TB1_IO_047;
  assign rx_pin[350] = mb1_FA2_TA2_IO_046_mb1_FB2_TB1_IO_044;
  assign rx_pin[351] = mb1_FA2_TA2_IO_047_mb1_FB2_TB1_IO_045;
  assign rx_pin[352] = mb1_FA2_TA2_IO_048_mb1_FB2_TB1_IO_062;
  assign rx_pin[353] = mb1_FA2_TA2_IO_049_mb1_FB2_TB1_IO_063;
  assign rx_pin[354] = mb1_FA2_TA2_IO_050_mb1_FB2_TB1_IO_040;
  assign rx_pin[355] = mb1_FA2_TA2_IO_051_mb1_FB2_TB1_IO_041;
  assign rx_pin[356] = mb1_FA2_TA2_IO_052_mb1_FB2_TB1_IO_038;
  assign rx_pin[357] = mb1_FA2_TA2_IO_053_mb1_FB2_TB1_IO_039;
  assign rx_pin[358] = mb1_FA2_TA2_IO_054_mb1_FB2_TB1_IO_056;
  assign rx_pin[359] = mb1_FA2_TA2_IO_055_mb1_FB2_TB1_IO_057;
  assign rx_pin[360] = mb1_FA2_TA2_IO_056_mb1_FB2_TB1_IO_054;
  assign rx_pin[361] = mb1_FA2_TA2_IO_057_mb1_FB2_TB1_IO_055;
  assign rx_pin[362] = mb1_FA2_TA2_IO_058_mb1_FB2_TB1_IO_072;
  assign rx_pin[363] = mb1_FA2_TA2_IO_059_mb1_FB2_TB1_IO_073;
  assign rx_pin[364] = mb1_FA2_TA2_IO_060_mb1_FB2_TB1_IO_070;
  assign rx_pin[365] = mb1_FA2_TA2_IO_061_mb1_FB2_TB1_IO_071;
  assign rx_pin[366] = mb1_FA2_TA2_IO_062_mb1_FB2_TB1_IO_048;
  assign rx_pin[367] = mb1_FA2_TA2_IO_063_mb1_FB2_TB1_IO_049;
  assign rx_pin[368] = mb1_FA2_TA2_IO_064_mb1_FB2_TB1_IO_066;
  assign rx_pin[369] = mb1_FA2_TA2_IO_065_mb1_FB2_TB1_IO_067;
  assign rx_pin[370] = mb1_FA2_TA2_IO_066_mb1_FB2_TB1_IO_064;
  assign rx_pin[371] = mb1_FA2_TA2_IO_067_mb1_FB2_TB1_IO_065;
  assign rx_pin[372] = mb1_FA2_TA2_IO_068_mb1_FB2_TB1_IO_082;
  assign rx_pin[373] = mb1_FA2_TA2_IO_069_mb1_FB2_TB1_IO_083;
  assign rx_pin[374] = mb1_FA2_TA2_IO_070_mb1_FB2_TB1_IO_060;
  assign rx_pin[375] = mb1_FA2_TA2_IO_071_mb1_FB2_TB1_IO_061;
  assign rx_pin[376] = mb1_FA2_TA2_IO_072_mb1_FB2_TB1_IO_058;
  assign rx_pin[377] = mb1_FA2_TA2_IO_073_mb1_FB2_TB1_IO_059;
  assign rx_pin[378] = mb1_FA2_TA2_IO_074_mb1_FB2_TB1_IO_076;
  assign rx_pin[379] = mb1_FA2_TA2_IO_075_mb1_FB2_TB1_IO_077;
  assign rx_pin[380] = mb1_FA2_TA2_IO_076_mb1_FB2_TB1_IO_074;
  assign rx_pin[381] = mb1_FA2_TA2_IO_077_mb1_FB2_TB1_IO_075;
  assign rx_pin[382] = mb1_FA2_TA2_IO_078_mb1_FB2_TB1_IO_092;
  assign rx_pin[383] = mb1_FA2_TA2_IO_079_mb1_FB2_TB1_IO_093;
  assign rx_pin[384] = mb1_FA2_TA2_IO_080_mb1_FB2_TB1_IO_090;
  assign rx_pin[385] = mb1_FA2_TA2_IO_081_mb1_FB2_TB1_IO_091;
  assign rx_pin[386] = mb1_FA2_TA2_IO_082_mb1_FB2_TB1_IO_068;
  assign rx_pin[387] = mb1_FA2_TA2_IO_083_mb1_FB2_TB1_IO_069;
  assign rx_pin[388] = mb1_FA2_TA2_IO_084_mb1_FB2_TB1_IO_086;
  assign rx_pin[389] = mb1_FA2_TA2_IO_085_mb1_FB2_TB1_IO_087;
  assign rx_pin[390] = mb1_FA2_TA2_IO_086_mb1_FB2_TB1_IO_084;
  assign rx_pin[391] = mb1_FA2_TA2_IO_087_mb1_FB2_TB1_IO_085;
  assign rx_pin[392] = mb1_FA2_TA2_IO_088_mb1_FB2_TB1_IO_102;
  assign rx_pin[393] = mb1_FA2_TA2_IO_089_mb1_FB2_TB1_IO_103;
  assign rx_pin[394] = mb1_FA2_TA2_IO_090_mb1_FB2_TB1_IO_080;
  assign rx_pin[395] = mb1_FA2_TA2_IO_091_mb1_FB2_TB1_IO_081;
  assign rx_pin[396] = mb1_FA2_TA2_IO_092_mb1_FB2_TB1_IO_078;
  assign rx_pin[397] = mb1_FA2_TA2_IO_093_mb1_FB2_TB1_IO_079;
  assign rx_pin[398] = mb1_FA2_TA2_IO_094_mb1_FB2_TB1_IO_096;
  assign rx_pin[399] = mb1_FA2_TA2_IO_095_mb1_FB2_TB1_IO_097;
  assign rx_pin[400] = mb1_FA2_TA2_IO_096_mb1_FB2_TB1_IO_094;
  assign rx_pin[401] = mb1_FA2_TA2_IO_097_mb1_FB2_TB1_IO_095;
  assign rx_pin[402] = mb1_FA2_TA2_IO_098_mb1_FB2_TB1_IO_112;
  assign rx_pin[403] = mb1_FA2_TA2_IO_099_mb1_FB2_TB1_IO_113;
  assign rx_pin[404] = mb1_FA2_TA2_IO_100_mb1_FB2_TB1_IO_110;
  assign rx_pin[405] = mb1_FA2_TA2_IO_101_mb1_FB2_TB1_IO_111;
  assign rx_pin[406] = mb1_FA2_TA2_IO_102_mb1_FB2_TB1_IO_088;
  assign rx_pin[407] = mb1_FA2_TA2_IO_103_mb1_FB2_TB1_IO_089;
  assign rx_pin[408] = mb1_FA2_TA2_IO_104_mb1_FB2_TB1_IO_106;
  assign rx_pin[409] = mb1_FA2_TA2_IO_105_mb1_FB2_TB1_IO_107;
  assign rx_pin[410] = mb1_FA2_TA2_IO_106_mb1_FB2_TB1_IO_104;
  assign rx_pin[411] = mb1_FA2_TA2_IO_107_mb1_FB2_TB1_IO_105;
  assign rx_pin[412] = mb1_FA2_TA2_IO_108_mb1_FB2_TB1_IO_122;
  assign rx_pin[413] = mb1_FA2_TA2_IO_109_mb1_FB2_TB1_IO_123;
  assign rx_pin[414] = mb1_FA2_TA2_IO_110_mb1_FB2_TB1_IO_100;
  assign rx_pin[415] = mb1_FA2_TA2_IO_111_mb1_FB2_TB1_IO_101;
  assign rx_pin[416] = mb1_FA2_TA2_IO_112_mb1_FB2_TB1_IO_098;
  assign rx_pin[417] = mb1_FA2_TA2_IO_113_mb1_FB2_TB1_IO_099;
  assign rx_pin[418] = mb1_FA2_TA2_IO_114_mb1_FB2_TB1_IO_116;
  assign rx_pin[419] = mb1_FA2_TA2_IO_115_mb1_FB2_TB1_IO_117;
  assign rx_pin[420] = mb1_FA2_TA2_IO_116_mb1_FB2_TB1_IO_114;
  assign rx_pin[421] = mb1_FA2_TA2_IO_117_mb1_FB2_TB1_IO_115;
  assign rx_pin[422] = mb1_FA2_TA2_IO_118_mb1_FB2_TB1_IO_132;
  assign rx_pin[423] = mb1_FA2_TA2_IO_119_mb1_FB2_TB1_IO_133;
  assign rx_pin[424] = mb1_FA2_TA2_IO_120_mb1_FB2_TB1_IO_130;
  assign rx_pin[425] = mb1_FA2_TA2_IO_121_mb1_FB2_TB1_IO_131;
  assign rx_pin[426] = mb1_FA2_TA2_IO_122_mb1_FB2_TB1_IO_108;
  assign rx_pin[427] = mb1_FA2_TA2_IO_123_mb1_FB2_TB1_IO_109;
  assign rx_pin[428] = mb1_FA2_TA2_IO_124_mb1_FB2_TB1_IO_126;
  assign rx_pin[429] = mb1_FA2_TA2_IO_125_mb1_FB2_TB1_IO_127;
  assign rx_pin[430] = mb1_FA2_TA2_IO_126_mb1_FB2_TB1_IO_124;
  assign rx_pin[431] = mb1_FA2_TA2_IO_127_mb1_FB2_TB1_IO_125;
  assign rx_pin[432] = mb1_FA2_TA2_IO_130_mb1_FB2_TB1_IO_120;
  assign rx_pin[433] = mb1_FA2_TA2_IO_131_mb1_FB2_TB1_IO_121;
  assign rx_pin[434] = mb1_FA2_TA2_IO_132_mb1_FB2_TB1_IO_118;
  assign rx_pin[435] = mb1_FA2_TA2_IO_133_mb1_FB2_TB1_IO_119;
  assign rx_pin[436] = mb1_FA2_TA2_IO_134_mb1_FB2_TB1_IO_136;
  assign rx_pin[437] = mb1_FA2_TA2_IO_136_mb1_FB2_TB1_IO_134;
  assign rx_pin[438] = mb1_FA2_TB2_CLKIO_N_0_mb1_FB2_TB2_CLKIO_N_7;
  assign rx_pin[439] = mb1_FA2_TB2_CLKIO_N_1_mb1_FB2_TB2_CLKIO_N_6;
  assign rx_pin[440] = mb1_FA2_TB2_CLKIO_N_2_mb1_FB2_TB2_CLKIO_N_4;
  assign rx_pin[441] = mb1_FA2_TB2_CLKIO_N_3_mb1_FB2_TB2_CLKIO_N_3;
  assign rx_pin[442] = mb1_FA2_TB2_CLKIO_N_4_mb1_FB2_TB2_CLKIO_N_2;
  assign rx_pin[443] = mb1_FA2_TB2_CLKIO_N_5_mb1_FB2_TB2_IO_010;
  assign rx_pin[444] = mb1_FA2_TB2_CLKIO_N_6_mb1_FB2_TB2_CLKIO_N_1;
  assign rx_pin[445] = mb1_FA2_TB2_CLKIO_N_7_mb1_FB2_TB2_CLKIO_N_0;
  assign rx_pin[446] = mb1_FA2_TB2_CLKIO_P_0_mb1_FB2_TB2_CLKIO_P_7;
  assign rx_pin[447] = mb1_FA2_TB2_CLKIO_P_1_mb1_FB2_TB2_CLKIO_P_6;
  assign rx_pin[448] = mb1_FA2_TB2_CLKIO_P_2_mb1_FB2_TB2_CLKIO_P_4;
  assign rx_pin[449] = mb1_FA2_TB2_CLKIO_P_3_mb1_FB2_TB2_CLKIO_P_3;
  assign rx_pin[450] = mb1_FA2_TB2_CLKIO_P_4_mb1_FB2_TB2_CLKIO_P_2;
  assign rx_pin[451] = mb1_FA2_TB2_CLKIO_P_5_mb1_FB2_TB2_IO_011;
  assign rx_pin[452] = mb1_FA2_TB2_CLKIO_P_6_mb1_FB2_TB2_CLKIO_P_1;
  assign rx_pin[453] = mb1_FA2_TB2_CLKIO_P_7_mb1_FB2_TB2_CLKIO_P_0;
  assign rx_pin[454] = mb1_FA2_TB2_IO_004_mb1_FB2_TB2_IO_006;
  assign rx_pin[455] = mb1_FA2_TB2_IO_005_mb1_FB2_TB2_IO_007;
  assign rx_pin[456] = mb1_FA2_TB2_IO_006_mb1_FB2_TB2_IO_004;
  assign rx_pin[457] = mb1_FA2_TB2_IO_007_mb1_FB2_TB2_IO_005;
  assign rx_pin[458] = mb1_FA2_TB2_IO_008_mb1_FB2_TB2_IO_022;
  assign rx_pin[459] = mb1_FA2_TB2_IO_009_mb1_FB2_TB2_IO_023;
  assign rx_pin[460] = mb1_FA2_TB2_IO_010_mb1_FB2_TB2_CLKIO_N_5;
  assign rx_pin[461] = mb1_FA2_TB2_IO_011_mb1_FB2_TB2_CLKIO_P_5;
  assign rx_pin[462] = mb1_FA2_TB2_IO_012_mb1_FB2_TB2_IO_012;
  assign rx_pin[463] = mb1_FA2_TB2_IO_013_mb1_FB2_TB2_IO_013;
  assign rx_pin[464] = mb1_FA2_TB2_IO_014_mb1_FB2_TB2_IO_016;
  assign rx_pin[465] = mb1_FA2_TB2_IO_015_mb1_FB2_TB2_IO_017;
  assign rx_pin[466] = mb1_FA2_TB2_IO_016_mb1_FB2_TB2_IO_014;
  assign rx_pin[467] = mb1_FA2_TB2_IO_017_mb1_FB2_TB2_IO_015;
  assign rx_pin[468] = mb1_FA2_TB2_IO_018_mb1_FB2_TB2_IO_032;
  assign rx_pin[469] = mb1_FA2_TB2_IO_019_mb1_FB2_TB2_IO_033;
  assign rx_pin[470] = mb1_FA2_TB2_IO_020_mb1_FB2_TB2_IO_030;
  assign rx_pin[471] = mb1_FA2_TB2_IO_021_mb1_FB2_TB2_IO_031;
  assign rx_pin[472] = mb1_FA2_TB2_IO_022_mb1_FB2_TB2_IO_008;
  assign rx_pin[473] = mb1_FA2_TB2_IO_023_mb1_FB2_TB2_IO_009;
  assign rx_pin[474] = mb1_FA2_TB2_IO_024_mb1_FB2_TB2_IO_026;
  assign rx_pin[475] = mb1_FA2_TB2_IO_025_mb1_FB2_TB2_IO_027;
  assign rx_pin[476] = mb1_FA2_TB2_IO_026_mb1_FB2_TB2_IO_024;
  assign rx_pin[477] = mb1_FA2_TB2_IO_027_mb1_FB2_TB2_IO_025;
  assign rx_pin[478] = mb1_FA2_TB2_IO_028_mb1_FB2_TB2_IO_042;
  assign rx_pin[479] = mb1_FA2_TB2_IO_029_mb1_FB2_TB2_IO_043;
  assign rx_pin[480] = mb1_FA2_TB2_IO_030_mb1_FB2_TB2_IO_020;
  assign rx_pin[481] = mb1_FA2_TB2_IO_031_mb1_FB2_TB2_IO_021;
  assign rx_pin[482] = mb1_FA2_TB2_IO_032_mb1_FB2_TB2_IO_018;
  assign rx_pin[483] = mb1_FA2_TB2_IO_033_mb1_FB2_TB2_IO_019;
  assign rx_pin[484] = mb1_FA2_TB2_IO_034_mb1_FB2_TB2_IO_036;
  assign rx_pin[485] = mb1_FA2_TB2_IO_035_mb1_FB2_TB2_IO_037;
  assign rx_pin[486] = mb1_FA2_TB2_IO_036_mb1_FB2_TB2_IO_034;
  assign rx_pin[487] = mb1_FA2_TB2_IO_037_mb1_FB2_TB2_IO_035;
  assign rx_pin[488] = mb1_FA2_TB2_IO_038_mb1_FB2_TB2_IO_052;
  assign rx_pin[489] = mb1_FA2_TB2_IO_039_mb1_FB2_TB2_IO_053;
  assign rx_pin[490] = mb1_FA2_TB2_IO_040_mb1_FB2_TB2_IO_050;
  assign rx_pin[491] = mb1_FA2_TB2_IO_041_mb1_FB2_TB2_IO_051;
  assign rx_pin[492] = mb1_FA2_TB2_IO_042_mb1_FB2_TB2_IO_028;
  assign rx_pin[493] = mb1_FA2_TB2_IO_043_mb1_FB2_TB2_IO_029;
  assign rx_pin[494] = mb1_FA2_TB2_IO_044_mb1_FB2_TB2_IO_046;
  assign rx_pin[495] = mb1_FA2_TB2_IO_045_mb1_FB2_TB2_IO_047;
  assign rx_pin[496] = mb1_FA2_TB2_IO_046_mb1_FB2_TB2_IO_044;
  assign rx_pin[497] = mb1_FA2_TB2_IO_047_mb1_FB2_TB2_IO_045;
  assign rx_pin[498] = mb1_FA2_TB2_IO_048_mb1_FB2_TB2_IO_062;
  assign rx_pin[499] = mb1_FA2_TB2_IO_049_mb1_FB2_TB2_IO_063;
  assign rx_pin[500] = mb1_FA2_TB2_IO_050_mb1_FB2_TB2_IO_040;
  assign rx_pin[501] = mb1_FA2_TB2_IO_051_mb1_FB2_TB2_IO_041;
  assign rx_pin[502] = mb1_FA2_TB2_IO_052_mb1_FB2_TB2_IO_038;
  assign rx_pin[503] = mb1_FA2_TB2_IO_053_mb1_FB2_TB2_IO_039;
  assign rx_pin[504] = mb1_FA2_TB2_IO_054_mb1_FB2_TB2_IO_056;
  assign rx_pin[505] = mb1_FA2_TB2_IO_055_mb1_FB2_TB2_IO_057;
  assign rx_pin[506] = mb1_FA2_TB2_IO_056_mb1_FB2_TB2_IO_054;
  assign rx_pin[507] = mb1_FA2_TB2_IO_057_mb1_FB2_TB2_IO_055;
  assign rx_pin[508] = mb1_FA2_TB2_IO_058_mb1_FB2_TB2_IO_072;
  assign rx_pin[509] = mb1_FA2_TB2_IO_059_mb1_FB2_TB2_IO_073;
  assign rx_pin[510] = mb1_FA2_TB2_IO_060_mb1_FB2_TB2_IO_070;
  assign rx_pin[511] = mb1_FA2_TB2_IO_061_mb1_FB2_TB2_IO_071;
  assign rx_pin[512] = mb1_FA2_TB2_IO_062_mb1_FB2_TB2_IO_048;
  assign rx_pin[513] = mb1_FA2_TB2_IO_063_mb1_FB2_TB2_IO_049;
  assign rx_pin[514] = mb1_FA2_TB2_IO_064_mb1_FB2_TB2_IO_066;
  assign rx_pin[515] = mb1_FA2_TB2_IO_065_mb1_FB2_TB2_IO_067;
  assign rx_pin[516] = mb1_FA2_TB2_IO_066_mb1_FB2_TB2_IO_064;
  assign rx_pin[517] = mb1_FA2_TB2_IO_067_mb1_FB2_TB2_IO_065;
  assign rx_pin[518] = mb1_FA2_TB2_IO_068_mb1_FB2_TB2_IO_082;
  assign rx_pin[519] = mb1_FA2_TB2_IO_069_mb1_FB2_TB2_IO_083;
  assign rx_pin[520] = mb1_FA2_TB2_IO_070_mb1_FB2_TB2_IO_060;
  assign rx_pin[521] = mb1_FA2_TB2_IO_071_mb1_FB2_TB2_IO_061;
  assign rx_pin[522] = mb1_FA2_TB2_IO_072_mb1_FB2_TB2_IO_058;
  assign rx_pin[523] = mb1_FA2_TB2_IO_073_mb1_FB2_TB2_IO_059;
  assign rx_pin[524] = mb1_FA2_TB2_IO_074_mb1_FB2_TB2_IO_076;
  assign rx_pin[525] = mb1_FA2_TB2_IO_075_mb1_FB2_TB2_IO_077;
  assign rx_pin[526] = mb1_FA2_TB2_IO_076_mb1_FB2_TB2_IO_074;
  assign rx_pin[527] = mb1_FA2_TB2_IO_077_mb1_FB2_TB2_IO_075;
  assign rx_pin[528] = mb1_FA2_TB2_IO_078_mb1_FB2_TB2_IO_092;
  assign rx_pin[529] = mb1_FA2_TB2_IO_079_mb1_FB2_TB2_IO_093;
  assign rx_pin[530] = mb1_FA2_TB2_IO_080_mb1_FB2_TB2_IO_090;
  assign rx_pin[531] = mb1_FA2_TB2_IO_081_mb1_FB2_TB2_IO_091;
  assign rx_pin[532] = mb1_FA2_TB2_IO_082_mb1_FB2_TB2_IO_068;
  assign rx_pin[533] = mb1_FA2_TB2_IO_083_mb1_FB2_TB2_IO_069;
  assign rx_pin[534] = mb1_FA2_TB2_IO_084_mb1_FB2_TB2_IO_086;
  assign rx_pin[535] = mb1_FA2_TB2_IO_085_mb1_FB2_TB2_IO_087;
  assign rx_pin[536] = mb1_FA2_TB2_IO_086_mb1_FB2_TB2_IO_084;
  assign rx_pin[537] = mb1_FA2_TB2_IO_087_mb1_FB2_TB2_IO_085;
  assign rx_pin[538] = mb1_FA2_TB2_IO_088_mb1_FB2_TB2_IO_102;
  assign rx_pin[539] = mb1_FA2_TB2_IO_089_mb1_FB2_TB2_IO_103;
  assign rx_pin[540] = mb1_FA2_TB2_IO_090_mb1_FB2_TB2_IO_080;
  assign rx_pin[541] = mb1_FA2_TB2_IO_091_mb1_FB2_TB2_IO_081;
  assign rx_pin[542] = mb1_FA2_TB2_IO_092_mb1_FB2_TB2_IO_078;
  assign rx_pin[543] = mb1_FA2_TB2_IO_093_mb1_FB2_TB2_IO_079;
  assign rx_pin[544] = mb1_FA2_TB2_IO_094_mb1_FB2_TB2_IO_096;
  assign rx_pin[545] = mb1_FA2_TB2_IO_095_mb1_FB2_TB2_IO_097;
  assign rx_pin[546] = mb1_FA2_TB2_IO_096_mb1_FB2_TB2_IO_094;
  assign rx_pin[547] = mb1_FA2_TB2_IO_097_mb1_FB2_TB2_IO_095;
  assign rx_pin[548] = mb1_FA2_TB2_IO_098_mb1_FB2_TB2_IO_112;
  assign rx_pin[549] = mb1_FA2_TB2_IO_099_mb1_FB2_TB2_IO_113;
  assign rx_pin[550] = mb1_FA2_TB2_IO_100_mb1_FB2_TB2_IO_110;
  assign rx_pin[551] = mb1_FA2_TB2_IO_101_mb1_FB2_TB2_IO_111;
  assign rx_pin[552] = mb1_FA2_TB2_IO_102_mb1_FB2_TB2_IO_088;
  assign rx_pin[553] = mb1_FA2_TB2_IO_103_mb1_FB2_TB2_IO_089;
  assign rx_pin[554] = mb1_FA2_TB2_IO_104_mb1_FB2_TB2_IO_106;
  assign rx_pin[555] = mb1_FA2_TB2_IO_105_mb1_FB2_TB2_IO_107;
  assign rx_pin[556] = mb1_FA2_TB2_IO_106_mb1_FB2_TB2_IO_104;
  assign rx_pin[557] = mb1_FA2_TB2_IO_107_mb1_FB2_TB2_IO_105;
  assign rx_pin[558] = mb1_FA2_TB2_IO_108_mb1_FB2_TB2_IO_122;
  assign rx_pin[559] = mb1_FA2_TB2_IO_109_mb1_FB2_TB2_IO_123;
  assign rx_pin[560] = mb1_FA2_TB2_IO_110_mb1_FB2_TB2_IO_100;
  assign rx_pin[561] = mb1_FA2_TB2_IO_111_mb1_FB2_TB2_IO_101;
  assign rx_pin[562] = mb1_FA2_TB2_IO_112_mb1_FB2_TB2_IO_098;
  assign rx_pin[563] = mb1_FA2_TB2_IO_113_mb1_FB2_TB2_IO_099;
  assign rx_pin[564] = mb1_FA2_TB2_IO_114_mb1_FB2_TB2_IO_116;
  assign rx_pin[565] = mb1_FA2_TB2_IO_115_mb1_FB2_TB2_IO_117;
  assign rx_pin[566] = mb1_FA2_TB2_IO_116_mb1_FB2_TB2_IO_114;
  assign rx_pin[567] = mb1_FA2_TB2_IO_117_mb1_FB2_TB2_IO_115;
  assign rx_pin[568] = mb1_FA2_TB2_IO_118_mb1_FB2_TB2_IO_132;
  assign rx_pin[569] = mb1_FA2_TB2_IO_119_mb1_FB2_TB2_IO_133;
  assign rx_pin[570] = mb1_FA2_TB2_IO_120_mb1_FB2_TB2_IO_130;
  assign rx_pin[571] = mb1_FA2_TB2_IO_121_mb1_FB2_TB2_IO_131;
  assign rx_pin[572] = mb1_FA2_TB2_IO_122_mb1_FB2_TB2_IO_108;
  assign rx_pin[573] = mb1_FA2_TB2_IO_123_mb1_FB2_TB2_IO_109;
  assign rx_pin[574] = mb1_FA2_TB2_IO_124_mb1_FB2_TB2_IO_126;
  assign rx_pin[575] = mb1_FA2_TB2_IO_125_mb1_FB2_TB2_IO_127;
  assign rx_pin[576] = mb1_FA2_TB2_IO_126_mb1_FB2_TB2_IO_124;
  assign rx_pin[577] = mb1_FA2_TB2_IO_127_mb1_FB2_TB2_IO_125;
  assign rx_pin[578] = mb1_FA2_TB2_IO_130_mb1_FB2_TB2_IO_120;
  assign rx_pin[579] = mb1_FA2_TB2_IO_131_mb1_FB2_TB2_IO_121;
  assign rx_pin[580] = mb1_FA2_TB2_IO_132_mb1_FB2_TB2_IO_118;
  assign rx_pin[581] = mb1_FA2_TB2_IO_133_mb1_FB2_TB2_IO_119;
  assign rx_pin[582] = mb1_FA2_TB2_IO_134_mb1_FB2_TB2_IO_136;
  assign rx_pin[583] = mb1_FA2_TB2_IO_136_mb1_FB2_TB2_IO_134;
  assign rx_pin[584] = mb1_FA2_TA1_CLKIO_N_0_mb1_FB2_BA0_CLKIO_N_7;
  assign rx_pin[585] = mb1_FA2_TA1_CLKIO_N_1_mb1_FB2_BA0_CLKIO_N_6;
  assign rx_pin[586] = mb1_FA2_TA1_CLKIO_N_2_mb1_FB2_BA0_CLKIO_N_4;
  assign rx_pin[587] = mb1_FA2_TA1_CLKIO_N_3_mb1_FB2_BA0_CLKIO_N_3;
  assign rx_pin[588] = mb1_FA2_TA1_CLKIO_N_4_mb1_FB2_BA0_CLKIO_N_2;
  assign rx_pin[589] = mb1_FA2_TA1_CLKIO_N_5_mb1_FB2_BA0_IO_010;
  assign rx_pin[590] = mb1_FA2_TA1_CLKIO_N_6_mb1_FB2_BA0_CLKIO_N_1;
  assign rx_pin[591] = mb1_FA2_TA1_CLKIO_N_7_mb1_FB2_BA0_CLKIO_N_0;
  assign rx_pin[592] = mb1_FA2_TA1_CLKIO_P_0_mb1_FB2_BA0_CLKIO_P_7;
  assign rx_pin[593] = mb1_FA2_TA1_CLKIO_P_1_mb1_FB2_BA0_CLKIO_P_6;
  assign rx_pin[594] = mb1_FA2_TA1_CLKIO_P_2_mb1_FB2_BA0_CLKIO_P_4;
  assign rx_pin[595] = mb1_FA2_TA1_CLKIO_P_3_mb1_FB2_BA0_CLKIO_P_3;
  assign rx_pin[596] = mb1_FA2_TA1_CLKIO_P_4_mb1_FB2_BA0_CLKIO_P_2;
  assign rx_pin[597] = mb1_FA2_TA1_CLKIO_P_5_mb1_FB2_BA0_IO_011;
  assign rx_pin[598] = mb1_FA2_TA1_CLKIO_P_6_mb1_FB2_BA0_CLKIO_P_1;
  assign rx_pin[599] = mb1_FA2_TA1_CLKIO_P_7_mb1_FB2_BA0_CLKIO_P_0;
  assign rx_pin[600] = mb1_FA2_TA1_IO_004_mb1_FB2_BA0_IO_006;
  assign rx_pin[601] = mb1_FA2_TA1_IO_005_mb1_FB2_BA0_IO_007;
  assign rx_pin[602] = mb1_FA2_TA1_IO_006_mb1_FB2_BA0_IO_004;
  assign rx_pin[603] = mb1_FA2_TA1_IO_007_mb1_FB2_BA0_IO_005;
  assign rx_pin[604] = mb1_FA2_TA1_IO_008_mb1_FB2_BA0_IO_022;
  assign rx_pin[605] = mb1_FA2_TA1_IO_009_mb1_FB2_BA0_IO_023;
  assign rx_pin[606] = mb1_FA2_TA1_IO_010_mb1_FB2_BA0_CLKIO_N_5;
  assign rx_pin[607] = mb1_FA2_TA1_IO_011_mb1_FB2_BA0_CLKIO_P_5;
  assign rx_pin[608] = mb1_FA2_TA1_IO_012_mb1_FB2_BA0_IO_012;
  assign rx_pin[609] = mb1_FA2_TA1_IO_013_mb1_FB2_BA0_IO_013;
  assign rx_pin[610] = mb1_FA2_TA1_IO_014_mb1_FB2_BA0_IO_016;
  assign rx_pin[611] = mb1_FA2_TA1_IO_015_mb1_FB2_BA0_IO_017;
  assign rx_pin[612] = mb1_FA2_TA1_IO_016_mb1_FB2_BA0_IO_014;
  assign rx_pin[613] = mb1_FA2_TA1_IO_017_mb1_FB2_BA0_IO_015;
  assign rx_pin[614] = mb1_FA2_TA1_IO_018_mb1_FB2_BA0_IO_032;
  assign rx_pin[615] = mb1_FA2_TA1_IO_019_mb1_FB2_BA0_IO_033;
  assign rx_pin[616] = mb1_FA2_TA1_IO_020_mb1_FB2_BA0_IO_030;
  assign rx_pin[617] = mb1_FA2_TA1_IO_021_mb1_FB2_BA0_IO_031;
  assign rx_pin[618] = mb1_FA2_TA1_IO_022_mb1_FB2_BA0_IO_008;
  assign rx_pin[619] = mb1_FA2_TA1_IO_023_mb1_FB2_BA0_IO_009;
  assign rx_pin[620] = mb1_FA2_TA1_IO_024_mb1_FB2_BA0_IO_026;
  assign rx_pin[621] = mb1_FA2_TA1_IO_025_mb1_FB2_BA0_IO_027;
  assign rx_pin[622] = mb1_FA2_TA1_IO_026_mb1_FB2_BA0_IO_024;
  assign rx_pin[623] = mb1_FA2_TA1_IO_027_mb1_FB2_BA0_IO_025;
  assign rx_pin[624] = mb1_FA2_TA1_IO_028_mb1_FB2_BA0_IO_042;
  assign rx_pin[625] = mb1_FA2_TA1_IO_029_mb1_FB2_BA0_IO_043;
  assign rx_pin[626] = mb1_FA2_TA1_IO_030_mb1_FB2_BA0_IO_020;
  assign rx_pin[627] = mb1_FA2_TA1_IO_031_mb1_FB2_BA0_IO_021;
  assign rx_pin[628] = mb1_FA2_TA1_IO_032_mb1_FB2_BA0_IO_018;
  assign rx_pin[629] = mb1_FA2_TA1_IO_033_mb1_FB2_BA0_IO_019;
  assign rx_pin[630] = mb1_FA2_TA1_IO_034_mb1_FB2_BA0_IO_036;
  assign rx_pin[631] = mb1_FA2_TA1_IO_035_mb1_FB2_BA0_IO_037;
  assign rx_pin[632] = mb1_FA2_TA1_IO_036_mb1_FB2_BA0_IO_034;
  assign rx_pin[633] = mb1_FA2_TA1_IO_037_mb1_FB2_BA0_IO_035;
  assign rx_pin[634] = mb1_FA2_TA1_IO_038_mb1_FB2_BA0_IO_052;
  assign rx_pin[635] = mb1_FA2_TA1_IO_039_mb1_FB2_BA0_IO_053;
  assign rx_pin[636] = mb1_FA2_TA1_IO_040_mb1_FB2_BA0_IO_050;
  assign rx_pin[637] = mb1_FA2_TA1_IO_041_mb1_FB2_BA0_IO_051;
  assign rx_pin[638] = mb1_FA2_TA1_IO_042_mb1_FB2_BA0_IO_028;
  assign rx_pin[639] = mb1_FA2_TA1_IO_043_mb1_FB2_BA0_IO_029;
  assign rx_pin[640] = mb1_FA2_TA1_IO_044_mb1_FB2_BA0_IO_046;
  assign rx_pin[641] = mb1_FA2_TA1_IO_045_mb1_FB2_BA0_IO_047;
  assign rx_pin[642] = mb1_FA2_TA1_IO_046_mb1_FB2_BA0_IO_044;
  assign rx_pin[643] = mb1_FA2_TA1_IO_047_mb1_FB2_BA0_IO_045;
  assign rx_pin[644] = mb1_FA2_TA1_IO_048_mb1_FB2_BA0_IO_062;
  assign rx_pin[645] = mb1_FA2_TA1_IO_049_mb1_FB2_BA0_IO_063;
  assign rx_pin[646] = mb1_FA2_TA1_IO_050_mb1_FB2_BA0_IO_040;
  assign rx_pin[647] = mb1_FA2_TA1_IO_051_mb1_FB2_BA0_IO_041;
  assign rx_pin[648] = mb1_FA2_TA1_IO_052_mb1_FB2_BA0_IO_038;
  assign rx_pin[649] = mb1_FA2_TA1_IO_053_mb1_FB2_BA0_IO_039;
  assign rx_pin[650] = mb1_FA2_TA1_IO_054_mb1_FB2_BA0_IO_056;
  assign rx_pin[651] = mb1_FA2_TA1_IO_055_mb1_FB2_BA0_IO_057;
  assign rx_pin[652] = mb1_FA2_TA1_IO_056_mb1_FB2_BA0_IO_054;
  assign rx_pin[653] = mb1_FA2_TA1_IO_057_mb1_FB2_BA0_IO_055;
  assign rx_pin[654] = mb1_FA2_TA1_IO_058_mb1_FB2_BA0_IO_072;
  assign rx_pin[655] = mb1_FA2_TA1_IO_059_mb1_FB2_BA0_IO_073;
  assign rx_pin[656] = mb1_FA2_TA1_IO_060_mb1_FB2_BA0_IO_070;
  assign rx_pin[657] = mb1_FA2_TA1_IO_061_mb1_FB2_BA0_IO_071;
  assign rx_pin[658] = mb1_FA2_TA1_IO_062_mb1_FB2_BA0_IO_048;
  assign rx_pin[659] = mb1_FA2_TA1_IO_063_mb1_FB2_BA0_IO_049;
  assign rx_pin[660] = mb1_FA2_TA1_IO_064_mb1_FB2_BA0_IO_066;
  assign rx_pin[661] = mb1_FA2_TA1_IO_065_mb1_FB2_BA0_IO_067;
  assign rx_pin[662] = mb1_FA2_TA1_IO_066_mb1_FB2_BA0_IO_064;
  assign rx_pin[663] = mb1_FA2_TA1_IO_067_mb1_FB2_BA0_IO_065;
  assign rx_pin[664] = mb1_FA2_TA1_IO_068_mb1_FB2_BA0_IO_082;
  assign rx_pin[665] = mb1_FA2_TA1_IO_069_mb1_FB2_BA0_IO_083;
  assign rx_pin[666] = mb1_FA2_TA1_IO_070_mb1_FB2_BA0_IO_060;
  assign rx_pin[667] = mb1_FA2_TA1_IO_071_mb1_FB2_BA0_IO_061;
  assign rx_pin[668] = mb1_FA2_TA1_IO_072_mb1_FB2_BA0_IO_058;
  assign rx_pin[669] = mb1_FA2_TA1_IO_073_mb1_FB2_BA0_IO_059;
  assign rx_pin[670] = mb1_FA2_TA1_IO_074_mb1_FB2_BA0_IO_076;
  assign rx_pin[671] = mb1_FA2_TA1_IO_075_mb1_FB2_BA0_IO_077;
  assign rx_pin[672] = mb1_FA2_TA1_IO_076_mb1_FB2_BA0_IO_074;
  assign rx_pin[673] = mb1_FA2_TA1_IO_077_mb1_FB2_BA0_IO_075;
  assign rx_pin[674] = mb1_FA2_TA1_IO_078_mb1_FB2_BA0_IO_092;
  assign rx_pin[675] = mb1_FA2_TA1_IO_079_mb1_FB2_BA0_IO_093;
  assign rx_pin[676] = mb1_FA2_TA1_IO_080_mb1_FB2_BA0_IO_090;
  assign rx_pin[677] = mb1_FA2_TA1_IO_081_mb1_FB2_BA0_IO_091;
  assign rx_pin[678] = mb1_FA2_TA1_IO_082_mb1_FB2_BA0_IO_068;
  assign rx_pin[679] = mb1_FA2_TA1_IO_083_mb1_FB2_BA0_IO_069;
  assign rx_pin[680] = mb1_FA2_TA1_IO_084_mb1_FB2_BA0_IO_086;
  assign rx_pin[681] = mb1_FA2_TA1_IO_085_mb1_FB2_BA0_IO_087;
  assign rx_pin[682] = mb1_FA2_TA1_IO_086_mb1_FB2_BA0_IO_084;
  assign rx_pin[683] = mb1_FA2_TA1_IO_087_mb1_FB2_BA0_IO_085;
  assign rx_pin[684] = mb1_FA2_TA1_IO_088_mb1_FB2_BA0_IO_102;
  assign rx_pin[685] = mb1_FA2_TA1_IO_089_mb1_FB2_BA0_IO_103;
  assign rx_pin[686] = mb1_FA2_TA1_IO_090_mb1_FB2_BA0_IO_080;
  assign rx_pin[687] = mb1_FA2_TA1_IO_091_mb1_FB2_BA0_IO_081;
  assign rx_pin[688] = mb1_FA2_TA1_IO_092_mb1_FB2_BA0_IO_078;
  assign rx_pin[689] = mb1_FA2_TA1_IO_093_mb1_FB2_BA0_IO_079;
  assign rx_pin[690] = mb1_FA2_TA1_IO_094_mb1_FB2_BA0_IO_096;
  assign rx_pin[691] = mb1_FA2_TA1_IO_095_mb1_FB2_BA0_IO_097;
  assign rx_pin[692] = mb1_FA2_TA1_IO_096_mb1_FB2_BA0_IO_094;
  assign rx_pin[693] = mb1_FA2_TA1_IO_097_mb1_FB2_BA0_IO_095;
  assign rx_pin[694] = mb1_FA2_TA1_IO_098_mb1_FB2_BA0_IO_112;
  assign rx_pin[695] = mb1_FA2_TA1_IO_099_mb1_FB2_BA0_IO_113;
  assign rx_pin[696] = mb1_FA2_TA1_IO_100_mb1_FB2_BA0_IO_110;
  assign rx_pin[697] = mb1_FA2_TA1_IO_101_mb1_FB2_BA0_IO_111;
  assign rx_pin[698] = mb1_FA2_TA1_IO_102_mb1_FB2_BA0_IO_088;
  assign rx_pin[699] = mb1_FA2_TA1_IO_103_mb1_FB2_BA0_IO_089;
  assign rx_pin[700] = mb1_FA2_TA1_IO_104_mb1_FB2_BA0_IO_106;
  assign rx_pin[701] = mb1_FA2_TA1_IO_105_mb1_FB2_BA0_IO_107;
  assign rx_pin[702] = mb1_FA2_TA1_IO_106_mb1_FB2_BA0_IO_104;
  assign rx_pin[703] = mb1_FA2_TA1_IO_107_mb1_FB2_BA0_IO_105;
  assign rx_pin[704] = mb1_FA2_TA1_IO_108_mb1_FB2_BA0_IO_122;
  assign rx_pin[705] = mb1_FA2_TA1_IO_109_mb1_FB2_BA0_IO_123;
  assign rx_pin[706] = mb1_FA2_TA1_IO_110_mb1_FB2_BA0_IO_100;
  assign rx_pin[707] = mb1_FA2_TA1_IO_111_mb1_FB2_BA0_IO_101;
  assign rx_pin[708] = mb1_FA2_TA1_IO_112_mb1_FB2_BA0_IO_098;
  assign rx_pin[709] = mb1_FA2_TA1_IO_113_mb1_FB2_BA0_IO_099;
  assign rx_pin[710] = mb1_FA2_TA1_IO_114_mb1_FB2_BA0_IO_116;
  assign rx_pin[711] = mb1_FA2_TA1_IO_115_mb1_FB2_BA0_IO_117;
  assign rx_pin[712] = mb1_FA2_TA1_IO_116_mb1_FB2_BA0_IO_114;
  assign rx_pin[713] = mb1_FA2_TA1_IO_117_mb1_FB2_BA0_IO_115;
  assign rx_pin[714] = mb1_FA2_TA1_IO_118_mb1_FB2_BA0_IO_132;
  assign rx_pin[715] = mb1_FA2_TA1_IO_119_mb1_FB2_BA0_IO_133;
  assign rx_pin[716] = mb1_FA2_TA1_IO_120_mb1_FB2_BA0_IO_130;
  assign rx_pin[717] = mb1_FA2_TA1_IO_121_mb1_FB2_BA0_IO_131;
  assign rx_pin[718] = mb1_FA2_TA1_IO_122_mb1_FB2_BA0_IO_108;
  assign rx_pin[719] = mb1_FA2_TA1_IO_123_mb1_FB2_BA0_IO_109;
  assign rx_pin[720] = mb1_FA2_TA1_IO_124_mb1_FB2_BA0_IO_126;
  assign rx_pin[721] = mb1_FA2_TA1_IO_125_mb1_FB2_BA0_IO_127;
  assign rx_pin[722] = mb1_FA2_TA1_IO_126_mb1_FB2_BA0_IO_124;
  assign rx_pin[723] = mb1_FA2_TA1_IO_127_mb1_FB2_BA0_IO_125;
  assign rx_pin[724] = mb1_FA2_TA1_IO_130_mb1_FB2_BA0_IO_120;
  assign rx_pin[725] = mb1_FA2_TA1_IO_131_mb1_FB2_BA0_IO_121;
  assign rx_pin[726] = mb1_FA2_TA1_IO_132_mb1_FB2_BA0_IO_118;
  assign rx_pin[727] = mb1_FA2_TA1_IO_133_mb1_FB2_BA0_IO_119;
  assign rx_pin[728] = mb1_FA2_TA1_IO_134_mb1_FB2_BA0_IO_136;
  assign rx_pin[729] = mb1_FA2_TA1_IO_136_mb1_FB2_BA0_IO_134;
  assign rx_pin[730] = mb1_FA2_BB0_CLKIO_N_0_mb1_FB2_BA1_CLKIO_N_7;
  assign rx_pin[731] = mb1_FA2_BB0_CLKIO_N_1_mb1_FB2_BA1_CLKIO_N_6;
  assign rx_pin[732] = mb1_FA2_BB0_CLKIO_N_2_mb1_FB2_BA1_CLKIO_N_4;
  assign rx_pin[733] = mb1_FA2_BB0_CLKIO_N_3_mb1_FB2_BA1_CLKIO_N_3;
  assign rx_pin[734] = mb1_FA2_BB0_CLKIO_N_4_mb1_FB2_BA1_CLKIO_N_2;
  assign rx_pin[735] = mb1_FA2_BB0_CLKIO_N_5_mb1_FB2_BA1_IO_010;
  assign rx_pin[736] = mb1_FA2_BB0_CLKIO_N_6_mb1_FB2_BA1_CLKIO_N_1;
  assign rx_pin[737] = mb1_FA2_BB0_CLKIO_N_7_mb1_FB2_BA1_CLKIO_N_0;
  assign rx_pin[738] = mb1_FA2_BB0_CLKIO_P_0_mb1_FB2_BA1_CLKIO_P_7;
  assign rx_pin[739] = mb1_FA2_BB0_CLKIO_P_1_mb1_FB2_BA1_CLKIO_P_6;
  assign rx_pin[740] = mb1_FA2_BB0_CLKIO_P_2_mb1_FB2_BA1_CLKIO_P_4;
  assign rx_pin[741] = mb1_FA2_BB0_CLKIO_P_3_mb1_FB2_BA1_CLKIO_P_3;
  assign rx_pin[742] = mb1_FA2_BB0_CLKIO_P_4_mb1_FB2_BA1_CLKIO_P_2;
  assign rx_pin[743] = mb1_FA2_BB0_CLKIO_P_5_mb1_FB2_BA1_IO_011;
  assign rx_pin[744] = mb1_FA2_BB0_CLKIO_P_6_mb1_FB2_BA1_CLKIO_P_1;
  assign rx_pin[745] = mb1_FA2_BB0_CLKIO_P_7_mb1_FB2_BA1_CLKIO_P_0;
  assign rx_pin[746] = mb1_FA2_BB0_IO_004_mb1_FB2_BA1_IO_006;
  assign rx_pin[747] = mb1_FA2_BB0_IO_005_mb1_FB2_BA1_IO_007;
  assign rx_pin[748] = mb1_FA2_BB0_IO_006_mb1_FB2_BA1_IO_004;
  assign rx_pin[749] = mb1_FA2_BB0_IO_007_mb1_FB2_BA1_IO_005;
  assign rx_pin[750] = mb1_FA2_BB0_IO_008_mb1_FB2_BA1_IO_022;
  assign rx_pin[751] = mb1_FA2_BB0_IO_009_mb1_FB2_BA1_IO_023;
  assign rx_pin[752] = mb1_FA2_BB0_IO_010_mb1_FB2_BA1_CLKIO_N_5;
  assign rx_pin[753] = mb1_FA2_BB0_IO_011_mb1_FB2_BA1_CLKIO_P_5;
  assign rx_pin[754] = mb1_FA2_BB0_IO_012_mb1_FB2_BA1_IO_012;
  assign rx_pin[755] = mb1_FA2_BB0_IO_013_mb1_FB2_BA1_IO_013;
  assign rx_pin[756] = mb1_FA2_BB0_IO_014_mb1_FB2_BA1_IO_016;
  assign rx_pin[757] = mb1_FA2_BB0_IO_015_mb1_FB2_BA1_IO_017;
  assign rx_pin[758] = mb1_FA2_BB0_IO_016_mb1_FB2_BA1_IO_014;
  assign rx_pin[759] = mb1_FA2_BB0_IO_017_mb1_FB2_BA1_IO_015;
  assign rx_pin[760] = mb1_FA2_BB0_IO_018_mb1_FB2_BA1_IO_032;
  assign rx_pin[761] = mb1_FA2_BB0_IO_019_mb1_FB2_BA1_IO_033;
  assign rx_pin[762] = mb1_FA2_BB0_IO_020_mb1_FB2_BA1_IO_030;
  assign rx_pin[763] = mb1_FA2_BB0_IO_021_mb1_FB2_BA1_IO_031;
  assign rx_pin[764] = mb1_FA2_BB0_IO_022_mb1_FB2_BA1_IO_008;
  assign rx_pin[765] = mb1_FA2_BB0_IO_023_mb1_FB2_BA1_IO_009;
  assign rx_pin[766] = mb1_FA2_BB0_IO_024_mb1_FB2_BA1_IO_026;
  assign rx_pin[767] = mb1_FA2_BB0_IO_025_mb1_FB2_BA1_IO_027;
  assign rx_pin[768] = mb1_FA2_BB0_IO_026_mb1_FB2_BA1_IO_024;
  assign rx_pin[769] = mb1_FA2_BB0_IO_027_mb1_FB2_BA1_IO_025;
  assign rx_pin[770] = mb1_FA2_BB0_IO_028_mb1_FB2_BA1_IO_042;
  assign rx_pin[771] = mb1_FA2_BB0_IO_029_mb1_FB2_BA1_IO_043;
  assign rx_pin[772] = mb1_FA2_BB0_IO_030_mb1_FB2_BA1_IO_020;
  assign rx_pin[773] = mb1_FA2_BB0_IO_031_mb1_FB2_BA1_IO_021;
  assign rx_pin[774] = mb1_FA2_BB0_IO_032_mb1_FB2_BA1_IO_018;
  assign rx_pin[775] = mb1_FA2_BB0_IO_033_mb1_FB2_BA1_IO_019;
  assign rx_pin[776] = mb1_FA2_BB0_IO_034_mb1_FB2_BA1_IO_036;
  assign rx_pin[777] = mb1_FA2_BB0_IO_035_mb1_FB2_BA1_IO_037;
  assign rx_pin[778] = mb1_FA2_BB0_IO_036_mb1_FB2_BA1_IO_034;
  assign rx_pin[779] = mb1_FA2_BB0_IO_037_mb1_FB2_BA1_IO_035;
  assign rx_pin[780] = mb1_FA2_BB0_IO_038_mb1_FB2_BA1_IO_052;
  assign rx_pin[781] = mb1_FA2_BB0_IO_039_mb1_FB2_BA1_IO_053;
  assign rx_pin[782] = mb1_FA2_BB0_IO_040_mb1_FB2_BA1_IO_050;
  assign rx_pin[783] = mb1_FA2_BB0_IO_041_mb1_FB2_BA1_IO_051;
  assign rx_pin[784] = mb1_FA2_BB0_IO_042_mb1_FB2_BA1_IO_028;
  assign rx_pin[785] = mb1_FA2_BB0_IO_043_mb1_FB2_BA1_IO_029;
  assign rx_pin[786] = mb1_FA2_BB0_IO_044_mb1_FB2_BA1_IO_046;
  assign rx_pin[787] = mb1_FA2_BB0_IO_045_mb1_FB2_BA1_IO_047;
  assign rx_pin[788] = mb1_FA2_BB0_IO_046_mb1_FB2_BA1_IO_044;
  assign rx_pin[789] = mb1_FA2_BB0_IO_047_mb1_FB2_BA1_IO_045;
  assign rx_pin[790] = mb1_FA2_BB0_IO_048_mb1_FB2_BA1_IO_062;
  assign rx_pin[791] = mb1_FA2_BB0_IO_049_mb1_FB2_BA1_IO_063;
  assign rx_pin[792] = mb1_FA2_BB0_IO_050_mb1_FB2_BA1_IO_040;
  assign rx_pin[793] = mb1_FA2_BB0_IO_051_mb1_FB2_BA1_IO_041;
  assign rx_pin[794] = mb1_FA2_BB0_IO_052_mb1_FB2_BA1_IO_038;
  assign rx_pin[795] = mb1_FA2_BB0_IO_053_mb1_FB2_BA1_IO_039;
  assign rx_pin[796] = mb1_FA2_BB0_IO_054_mb1_FB2_BA1_IO_056;
  assign rx_pin[797] = mb1_FA2_BB0_IO_055_mb1_FB2_BA1_IO_057;
  assign rx_pin[798] = mb1_FA2_BB0_IO_056_mb1_FB2_BA1_IO_054;
  assign rx_pin[799] = mb1_FA2_BB0_IO_057_mb1_FB2_BA1_IO_055;
  assign rx_pin[800] = mb1_FA2_BB0_IO_058_mb1_FB2_BA1_IO_072;
  assign rx_pin[801] = mb1_FA2_BB0_IO_059_mb1_FB2_BA1_IO_073;
  assign rx_pin[802] = mb1_FA2_BB0_IO_060_mb1_FB2_BA1_IO_070;
  assign rx_pin[803] = mb1_FA2_BB0_IO_061_mb1_FB2_BA1_IO_071;
  assign rx_pin[804] = mb1_FA2_BB0_IO_062_mb1_FB2_BA1_IO_048;
  assign rx_pin[805] = mb1_FA2_BB0_IO_063_mb1_FB2_BA1_IO_049;
  assign rx_pin[806] = mb1_FA2_BB0_IO_064_mb1_FB2_BA1_IO_066;
  assign rx_pin[807] = mb1_FA2_BB0_IO_065_mb1_FB2_BA1_IO_067;
  assign rx_pin[808] = mb1_FA2_BB0_IO_066_mb1_FB2_BA1_IO_064;
  assign rx_pin[809] = mb1_FA2_BB0_IO_067_mb1_FB2_BA1_IO_065;
  assign rx_pin[810] = mb1_FA2_BB0_IO_068_mb1_FB2_BA1_IO_082;
  assign rx_pin[811] = mb1_FA2_BB0_IO_069_mb1_FB2_BA1_IO_083;
  assign rx_pin[812] = mb1_FA2_BB0_IO_070_mb1_FB2_BA1_IO_060;
  assign rx_pin[813] = mb1_FA2_BB0_IO_071_mb1_FB2_BA1_IO_061;
  assign rx_pin[814] = mb1_FA2_BB0_IO_072_mb1_FB2_BA1_IO_058;
  assign rx_pin[815] = mb1_FA2_BB0_IO_073_mb1_FB2_BA1_IO_059;
  assign rx_pin[816] = mb1_FA2_BB0_IO_074_mb1_FB2_BA1_IO_076;
  assign rx_pin[817] = mb1_FA2_BB0_IO_075_mb1_FB2_BA1_IO_077;
  assign rx_pin[818] = mb1_FA2_BB0_IO_076_mb1_FB2_BA1_IO_074;
  assign rx_pin[819] = mb1_FA2_BB0_IO_077_mb1_FB2_BA1_IO_075;
  assign rx_pin[820] = mb1_FA2_BB0_IO_078_mb1_FB2_BA1_IO_092;
  assign rx_pin[821] = mb1_FA2_BB0_IO_079_mb1_FB2_BA1_IO_093;
  assign rx_pin[822] = mb1_FA2_BB0_IO_080_mb1_FB2_BA1_IO_090;
  assign rx_pin[823] = mb1_FA2_BB0_IO_081_mb1_FB2_BA1_IO_091;
  assign rx_pin[824] = mb1_FA2_BB0_IO_082_mb1_FB2_BA1_IO_068;
  assign rx_pin[825] = mb1_FA2_BB0_IO_083_mb1_FB2_BA1_IO_069;
  assign rx_pin[826] = mb1_FA2_BB0_IO_084_mb1_FB2_BA1_IO_086;
  assign rx_pin[827] = mb1_FA2_BB0_IO_085_mb1_FB2_BA1_IO_087;
  assign rx_pin[828] = mb1_FA2_BB0_IO_086_mb1_FB2_BA1_IO_084;
  assign rx_pin[829] = mb1_FA2_BB0_IO_087_mb1_FB2_BA1_IO_085;
  assign rx_pin[830] = mb1_FA2_BB0_IO_088_mb1_FB2_BA1_IO_102;
  assign rx_pin[831] = mb1_FA2_BB0_IO_089_mb1_FB2_BA1_IO_103;
  assign rx_pin[832] = mb1_FA2_BB0_IO_090_mb1_FB2_BA1_IO_080;
  assign rx_pin[833] = mb1_FA2_BB0_IO_091_mb1_FB2_BA1_IO_081;
  assign rx_pin[834] = mb1_FA2_BB0_IO_092_mb1_FB2_BA1_IO_078;
  assign rx_pin[835] = mb1_FA2_BB0_IO_093_mb1_FB2_BA1_IO_079;
  assign rx_pin[836] = mb1_FA2_BB0_IO_094_mb1_FB2_BA1_IO_096;
  assign rx_pin[837] = mb1_FA2_BB0_IO_095_mb1_FB2_BA1_IO_097;
  assign rx_pin[838] = mb1_FA2_BB0_IO_096_mb1_FB2_BA1_IO_094;
  assign rx_pin[839] = mb1_FA2_BB0_IO_097_mb1_FB2_BA1_IO_095;
  assign rx_pin[840] = mb1_FA2_BB0_IO_098_mb1_FB2_BA1_IO_112;
  assign rx_pin[841] = mb1_FA2_BB0_IO_099_mb1_FB2_BA1_IO_113;
  assign rx_pin[842] = mb1_FA2_BB0_IO_100_mb1_FB2_BA1_IO_110;
  assign rx_pin[843] = mb1_FA2_BB0_IO_101_mb1_FB2_BA1_IO_111;
  assign rx_pin[844] = mb1_FA2_BB0_IO_102_mb1_FB2_BA1_IO_088;
  assign rx_pin[845] = mb1_FA2_BB0_IO_103_mb1_FB2_BA1_IO_089;
  assign rx_pin[846] = mb1_FA2_BB0_IO_104_mb1_FB2_BA1_IO_106;
  assign rx_pin[847] = mb1_FA2_BB0_IO_105_mb1_FB2_BA1_IO_107;
  assign rx_pin[848] = mb1_FA2_BB0_IO_106_mb1_FB2_BA1_IO_104;
  assign rx_pin[849] = mb1_FA2_BB0_IO_107_mb1_FB2_BA1_IO_105;
  assign rx_pin[850] = mb1_FA2_BB0_IO_108_mb1_FB2_BA1_IO_122;
  assign rx_pin[851] = mb1_FA2_BB0_IO_109_mb1_FB2_BA1_IO_123;
  assign rx_pin[852] = mb1_FA2_BB0_IO_110_mb1_FB2_BA1_IO_100;
  assign rx_pin[853] = mb1_FA2_BB0_IO_111_mb1_FB2_BA1_IO_101;
  assign rx_pin[854] = mb1_FA2_BB0_IO_112_mb1_FB2_BA1_IO_098;
  assign rx_pin[855] = mb1_FA2_BB0_IO_113_mb1_FB2_BA1_IO_099;
  assign rx_pin[856] = mb1_FA2_BB0_IO_114_mb1_FB2_BA1_IO_116;
  assign rx_pin[857] = mb1_FA2_BB0_IO_115_mb1_FB2_BA1_IO_117;
  assign rx_pin[858] = mb1_FA2_BB0_IO_116_mb1_FB2_BA1_IO_114;
  assign rx_pin[859] = mb1_FA2_BB0_IO_117_mb1_FB2_BA1_IO_115;
  assign rx_pin[860] = mb1_FA2_BB0_IO_118_mb1_FB2_BA1_IO_132;
  assign rx_pin[861] = mb1_FA2_BB0_IO_119_mb1_FB2_BA1_IO_133;
  assign rx_pin[862] = mb1_FA2_BB0_IO_120_mb1_FB2_BA1_IO_130;
  assign rx_pin[863] = mb1_FA2_BB0_IO_121_mb1_FB2_BA1_IO_131;
  assign rx_pin[864] = mb1_FA2_BB0_IO_122_mb1_FB2_BA1_IO_108;
  assign rx_pin[865] = mb1_FA2_BB0_IO_123_mb1_FB2_BA1_IO_109;
  assign rx_pin[866] = mb1_FA2_BB0_IO_124_mb1_FB2_BA1_IO_126;
  assign rx_pin[867] = mb1_FA2_BB0_IO_125_mb1_FB2_BA1_IO_127;
  assign rx_pin[868] = mb1_FA2_BB0_IO_126_mb1_FB2_BA1_IO_124;
  assign rx_pin[869] = mb1_FA2_BB0_IO_127_mb1_FB2_BA1_IO_125;
  assign rx_pin[870] = mb1_FA2_BB0_IO_130_mb1_FB2_BA1_IO_120;
  assign rx_pin[871] = mb1_FA2_BB0_IO_131_mb1_FB2_BA1_IO_121;
  assign rx_pin[872] = mb1_FA2_BB0_IO_132_mb1_FB2_BA1_IO_118;
  assign rx_pin[873] = mb1_FA2_BB0_IO_133_mb1_FB2_BA1_IO_119;
  assign rx_pin[874] = mb1_FA2_BB0_IO_134_mb1_FB2_BA1_IO_136;
  assign rx_pin[875] = mb1_FA2_BB0_IO_136_mb1_FB2_BA1_IO_134;
  assign rx_pin[876] = mb1_FA2_BA2_CLKIO_N_0_mb1_FB2_BA2_CLKIO_N_7;
  assign rx_pin[877] = mb1_FA2_BA2_CLKIO_N_1_mb1_FB2_BA2_CLKIO_N_6;
  assign rx_pin[878] = mb1_FA2_BA2_CLKIO_N_2_mb1_FB2_BA2_CLKIO_N_4;
  assign rx_pin[879] = mb1_FA2_BA2_CLKIO_N_3_mb1_FB2_BA2_CLKIO_N_3;
  assign rx_pin[880] = mb1_FA2_BA2_CLKIO_N_4_mb1_FB2_BA2_CLKIO_N_2;
  assign rx_pin[881] = mb1_FA2_BA2_CLKIO_N_5_mb1_FB2_BA2_IO_010;
  assign rx_pin[882] = mb1_FA2_BA2_CLKIO_N_6_mb1_FB2_BA2_CLKIO_N_1;
  assign rx_pin[883] = mb1_FA2_BA2_CLKIO_N_7_mb1_FB2_BA2_CLKIO_N_0;
  assign rx_pin[884] = mb1_FA2_BA2_CLKIO_P_0_mb1_FB2_BA2_CLKIO_P_7;
  assign rx_pin[885] = mb1_FA2_BA2_CLKIO_P_1_mb1_FB2_BA2_CLKIO_P_6;
  assign rx_pin[886] = mb1_FA2_BA2_CLKIO_P_2_mb1_FB2_BA2_CLKIO_P_4;
  assign rx_pin[887] = mb1_FA2_BA2_CLKIO_P_3_mb1_FB2_BA2_CLKIO_P_3;
  assign rx_pin[888] = mb1_FA2_BA2_CLKIO_P_4_mb1_FB2_BA2_CLKIO_P_2;
  assign rx_pin[889] = mb1_FA2_BA2_CLKIO_P_5_mb1_FB2_BA2_IO_011;
  assign rx_pin[890] = mb1_FA2_BA2_CLKIO_P_6_mb1_FB2_BA2_CLKIO_P_1;
  assign rx_pin[891] = mb1_FA2_BA2_CLKIO_P_7_mb1_FB2_BA2_CLKIO_P_0;
  assign rx_pin[892] = mb1_FA2_BA2_IO_004_mb1_FB2_BA2_IO_006;
  assign rx_pin[893] = mb1_FA2_BA2_IO_005_mb1_FB2_BA2_IO_007;
  assign rx_pin[894] = mb1_FA2_BA2_IO_006_mb1_FB2_BA2_IO_004;
  assign rx_pin[895] = mb1_FA2_BA2_IO_007_mb1_FB2_BA2_IO_005;
  assign rx_pin[896] = mb1_FA2_BA2_IO_008_mb1_FB2_BA2_IO_022;
  assign rx_pin[897] = mb1_FA2_BA2_IO_009_mb1_FB2_BA2_IO_023;
  assign rx_pin[898] = mb1_FA2_BA2_IO_010_mb1_FB2_BA2_CLKIO_N_5;
  assign rx_pin[899] = mb1_FA2_BA2_IO_011_mb1_FB2_BA2_CLKIO_P_5;
  assign rx_pin[900] = mb1_FA2_BA2_IO_012_mb1_FB2_BA2_IO_012;
  assign rx_pin[901] = mb1_FA2_BA2_IO_013_mb1_FB2_BA2_IO_013;
  assign rx_pin[902] = mb1_FA2_BA2_IO_014_mb1_FB2_BA2_IO_016;
  assign rx_pin[903] = mb1_FA2_BA2_IO_015_mb1_FB2_BA2_IO_017;
  assign rx_pin[904] = mb1_FA2_BA2_IO_016_mb1_FB2_BA2_IO_014;
  assign rx_pin[905] = mb1_FA2_BA2_IO_017_mb1_FB2_BA2_IO_015;
  assign rx_pin[906] = mb1_FA2_BA2_IO_018_mb1_FB2_BA2_IO_032;
  assign rx_pin[907] = mb1_FA2_BA2_IO_019_mb1_FB2_BA2_IO_033;
  assign rx_pin[908] = mb1_FA2_BA2_IO_020_mb1_FB2_BA2_IO_030;
  assign rx_pin[909] = mb1_FA2_BA2_IO_021_mb1_FB2_BA2_IO_031;
  assign rx_pin[910] = mb1_FA2_BA2_IO_022_mb1_FB2_BA2_IO_008;
  assign rx_pin[911] = mb1_FA2_BA2_IO_023_mb1_FB2_BA2_IO_009;
  assign rx_pin[912] = mb1_FA2_BA2_IO_024_mb1_FB2_BA2_IO_026;
  assign rx_pin[913] = mb1_FA2_BA2_IO_025_mb1_FB2_BA2_IO_027;
  assign rx_pin[914] = mb1_FA2_BA2_IO_026_mb1_FB2_BA2_IO_024;
  assign rx_pin[915] = mb1_FA2_BA2_IO_027_mb1_FB2_BA2_IO_025;
  assign rx_pin[916] = mb1_FA2_BA2_IO_028_mb1_FB2_BA2_IO_042;
  assign rx_pin[917] = mb1_FA2_BA2_IO_029_mb1_FB2_BA2_IO_043;
  assign rx_pin[918] = mb1_FA2_BA2_IO_030_mb1_FB2_BA2_IO_020;
  assign rx_pin[919] = mb1_FA2_BA2_IO_031_mb1_FB2_BA2_IO_021;
  assign rx_pin[920] = mb1_FA2_BA2_IO_032_mb1_FB2_BA2_IO_018;
  assign rx_pin[921] = mb1_FA2_BA2_IO_033_mb1_FB2_BA2_IO_019;
  assign rx_pin[922] = mb1_FA2_BA2_IO_034_mb1_FB2_BA2_IO_036;
  assign rx_pin[923] = mb1_FA2_BA2_IO_035_mb1_FB2_BA2_IO_037;
  assign rx_pin[924] = mb1_FA2_BA2_IO_036_mb1_FB2_BA2_IO_034;
  assign rx_pin[925] = mb1_FA2_BA2_IO_037_mb1_FB2_BA2_IO_035;
  assign rx_pin[926] = mb1_FA2_BA2_IO_038_mb1_FB2_BA2_IO_052;
  assign rx_pin[927] = mb1_FA2_BA2_IO_039_mb1_FB2_BA2_IO_053;
  assign rx_pin[928] = mb1_FA2_BA2_IO_040_mb1_FB2_BA2_IO_050;
  assign rx_pin[929] = mb1_FA2_BA2_IO_041_mb1_FB2_BA2_IO_051;
  assign rx_pin[930] = mb1_FA2_BA2_IO_042_mb1_FB2_BA2_IO_028;
  assign rx_pin[931] = mb1_FA2_BA2_IO_043_mb1_FB2_BA2_IO_029;
  assign rx_pin[932] = mb1_FA2_BA2_IO_044_mb1_FB2_BA2_IO_046;
  assign rx_pin[933] = mb1_FA2_BA2_IO_045_mb1_FB2_BA2_IO_047;
  assign rx_pin[934] = mb1_FA2_BA2_IO_046_mb1_FB2_BA2_IO_044;
  assign rx_pin[935] = mb1_FA2_BA2_IO_047_mb1_FB2_BA2_IO_045;
  assign rx_pin[936] = mb1_FA2_BA2_IO_048_mb1_FB2_BA2_IO_062;
  assign rx_pin[937] = mb1_FA2_BA2_IO_049_mb1_FB2_BA2_IO_063;
  assign rx_pin[938] = mb1_FA2_BA2_IO_050_mb1_FB2_BA2_IO_040;
  assign rx_pin[939] = mb1_FA2_BA2_IO_051_mb1_FB2_BA2_IO_041;
  assign rx_pin[940] = mb1_FA2_BA2_IO_052_mb1_FB2_BA2_IO_038;
  assign rx_pin[941] = mb1_FA2_BA2_IO_053_mb1_FB2_BA2_IO_039;
  assign rx_pin[942] = mb1_FA2_BA2_IO_054_mb1_FB2_BA2_IO_056;
  assign rx_pin[943] = mb1_FA2_BA2_IO_055_mb1_FB2_BA2_IO_057;
  assign rx_pin[944] = mb1_FA2_BA2_IO_056_mb1_FB2_BA2_IO_054;
  assign rx_pin[945] = mb1_FA2_BA2_IO_057_mb1_FB2_BA2_IO_055;
  assign rx_pin[946] = mb1_FA2_BA2_IO_058_mb1_FB2_BA2_IO_072;
  assign rx_pin[947] = mb1_FA2_BA2_IO_059_mb1_FB2_BA2_IO_073;
  assign rx_pin[948] = mb1_FA2_BA2_IO_060_mb1_FB2_BA2_IO_070;
  assign rx_pin[949] = mb1_FA2_BA2_IO_061_mb1_FB2_BA2_IO_071;
  assign rx_pin[950] = mb1_FA2_BA2_IO_062_mb1_FB2_BA2_IO_048;
  assign rx_pin[951] = mb1_FA2_BA2_IO_063_mb1_FB2_BA2_IO_049;
  assign rx_pin[952] = mb1_FA2_BA2_IO_064_mb1_FB2_BA2_IO_066;
  assign rx_pin[953] = mb1_FA2_BA2_IO_065_mb1_FB2_BA2_IO_067;
  assign rx_pin[954] = mb1_FA2_BA2_IO_066_mb1_FB2_BA2_IO_064;
  assign rx_pin[955] = mb1_FA2_BA2_IO_067_mb1_FB2_BA2_IO_065;
  assign rx_pin[956] = mb1_FA2_BA2_IO_068_mb1_FB2_BA2_IO_082;
  assign rx_pin[957] = mb1_FA2_BA2_IO_069_mb1_FB2_BA2_IO_083;
  assign rx_pin[958] = mb1_FA2_BA2_IO_070_mb1_FB2_BA2_IO_060;
  assign rx_pin[959] = mb1_FA2_BA2_IO_071_mb1_FB2_BA2_IO_061;
  assign rx_pin[960] = mb1_FA2_BA2_IO_072_mb1_FB2_BA2_IO_058;
  assign rx_pin[961] = mb1_FA2_BA2_IO_073_mb1_FB2_BA2_IO_059;
  assign rx_pin[962] = mb1_FA2_BA2_IO_074_mb1_FB2_BA2_IO_076;
  assign rx_pin[963] = mb1_FA2_BA2_IO_075_mb1_FB2_BA2_IO_077;
  assign rx_pin[964] = mb1_FA2_BA2_IO_076_mb1_FB2_BA2_IO_074;
  assign rx_pin[965] = mb1_FA2_BA2_IO_077_mb1_FB2_BA2_IO_075;
  assign rx_pin[966] = mb1_FA2_BA2_IO_078_mb1_FB2_BA2_IO_092;
  assign rx_pin[967] = mb1_FA2_BA2_IO_079_mb1_FB2_BA2_IO_093;
  assign rx_pin[968] = mb1_FA2_BA2_IO_080_mb1_FB2_BA2_IO_090;
  assign rx_pin[969] = mb1_FA2_BA2_IO_081_mb1_FB2_BA2_IO_091;
  assign rx_pin[970] = mb1_FA2_BA2_IO_082_mb1_FB2_BA2_IO_068;
  assign rx_pin[971] = mb1_FA2_BA2_IO_083_mb1_FB2_BA2_IO_069;
  assign rx_pin[972] = mb1_FA2_BA2_IO_084_mb1_FB2_BA2_IO_086;
  assign rx_pin[973] = mb1_FA2_BA2_IO_085_mb1_FB2_BA2_IO_087;
  assign rx_pin[974] = mb1_FA2_BA2_IO_086_mb1_FB2_BA2_IO_084;
  assign rx_pin[975] = mb1_FA2_BA2_IO_087_mb1_FB2_BA2_IO_085;
  assign rx_pin[976] = mb1_FA2_BA2_IO_088_mb1_FB2_BA2_IO_102;
  assign rx_pin[977] = mb1_FA2_BA2_IO_089_mb1_FB2_BA2_IO_103;
  assign rx_pin[978] = mb1_FA2_BA2_IO_090_mb1_FB2_BA2_IO_080;
  assign rx_pin[979] = mb1_FA2_BA2_IO_091_mb1_FB2_BA2_IO_081;
  assign rx_pin[980] = mb1_FA2_BA2_IO_092_mb1_FB2_BA2_IO_078;
  assign rx_pin[981] = mb1_FA2_BA2_IO_093_mb1_FB2_BA2_IO_079;
  assign rx_pin[982] = mb1_FA2_BA2_IO_094_mb1_FB2_BA2_IO_096;
  assign rx_pin[983] = mb1_FA2_BA2_IO_095_mb1_FB2_BA2_IO_097;
  assign rx_pin[984] = mb1_FA2_BA2_IO_096_mb1_FB2_BA2_IO_094;
  assign rx_pin[985] = mb1_FA2_BA2_IO_097_mb1_FB2_BA2_IO_095;
  assign rx_pin[986] = mb1_FA2_BA2_IO_098_mb1_FB2_BA2_IO_112;
  assign rx_pin[987] = mb1_FA2_BA2_IO_099_mb1_FB2_BA2_IO_113;
  assign rx_pin[988] = mb1_FA2_BA2_IO_100_mb1_FB2_BA2_IO_110;
  assign rx_pin[989] = mb1_FA2_BA2_IO_101_mb1_FB2_BA2_IO_111;
  assign rx_pin[990] = mb1_FA2_BA2_IO_102_mb1_FB2_BA2_IO_088;
  assign rx_pin[991] = mb1_FA2_BA2_IO_103_mb1_FB2_BA2_IO_089;
  assign rx_pin[992] = mb1_FA2_BA2_IO_104_mb1_FB2_BA2_IO_106;
  assign rx_pin[993] = mb1_FA2_BA2_IO_105_mb1_FB2_BA2_IO_107;
  assign rx_pin[994] = mb1_FA2_BA2_IO_106_mb1_FB2_BA2_IO_104;
  assign rx_pin[995] = mb1_FA2_BA2_IO_107_mb1_FB2_BA2_IO_105;
  assign rx_pin[996] = mb1_FA2_BA2_IO_108_mb1_FB2_BA2_IO_122;
  assign rx_pin[997] = mb1_FA2_BA2_IO_109_mb1_FB2_BA2_IO_123;
  assign rx_pin[998] = mb1_FA2_BA2_IO_110_mb1_FB2_BA2_IO_100;
  assign rx_pin[999] = mb1_FA2_BA2_IO_111_mb1_FB2_BA2_IO_101;
  assign rx_pin[1000] = mb1_FA2_BA2_IO_112_mb1_FB2_BA2_IO_098;
  assign rx_pin[1001] = mb1_FA2_BA2_IO_113_mb1_FB2_BA2_IO_099;
  assign rx_pin[1002] = mb1_FA2_BA2_IO_114_mb1_FB2_BA2_IO_116;
  assign rx_pin[1003] = mb1_FA2_BA2_IO_115_mb1_FB2_BA2_IO_117;
  assign rx_pin[1004] = mb1_FA2_BA2_IO_116_mb1_FB2_BA2_IO_114;
  assign rx_pin[1005] = mb1_FA2_BA2_IO_117_mb1_FB2_BA2_IO_115;
  assign rx_pin[1006] = mb1_FA2_BA2_IO_118_mb1_FB2_BA2_IO_132;
  assign rx_pin[1007] = mb1_FA2_BA2_IO_119_mb1_FB2_BA2_IO_133;
  assign rx_pin[1008] = mb1_FA2_BA2_IO_120_mb1_FB2_BA2_IO_130;
  assign rx_pin[1009] = mb1_FA2_BA2_IO_121_mb1_FB2_BA2_IO_131;
  assign rx_pin[1010] = mb1_FA2_BA2_IO_122_mb1_FB2_BA2_IO_108;
  assign rx_pin[1011] = mb1_FA2_BA2_IO_123_mb1_FB2_BA2_IO_109;
  assign rx_pin[1012] = mb1_FA2_BA2_IO_124_mb1_FB2_BA2_IO_126;
  assign rx_pin[1013] = mb1_FA2_BA2_IO_125_mb1_FB2_BA2_IO_127;
  assign rx_pin[1014] = mb1_FA2_BA2_IO_126_mb1_FB2_BA2_IO_124;
  assign rx_pin[1015] = mb1_FA2_BA2_IO_127_mb1_FB2_BA2_IO_125;
  assign rx_pin[1016] = mb1_FA2_BA2_IO_130_mb1_FB2_BA2_IO_120;
  assign rx_pin[1017] = mb1_FA2_BA2_IO_131_mb1_FB2_BA2_IO_121;
  assign rx_pin[1018] = mb1_FA2_BA2_IO_132_mb1_FB2_BA2_IO_118;
  assign rx_pin[1019] = mb1_FA2_BA2_IO_133_mb1_FB2_BA2_IO_119;
  assign rx_pin[1020] = mb1_FA2_BA2_IO_134_mb1_FB2_BA2_IO_136;
  assign rx_pin[1021] = mb1_FA2_BA2_IO_136_mb1_FB2_BA2_IO_134;
  assign rx_pin[1022] = mb1_FB1_TA1_CLKIO_N_0_mb1_FB2_BB0_CLKIO_N_7;
  assign rx_pin[1023] = mb1_FB1_TA1_CLKIO_N_1_mb1_FB2_BB0_CLKIO_N_6;
  assign rx_pin[1024] = mb1_FB1_TA1_CLKIO_N_2_mb1_FB2_BB0_CLKIO_N_4;
  assign rx_pin[1025] = mb1_FB1_TA1_CLKIO_N_3_mb1_FB2_BB0_CLKIO_N_3;
  assign rx_pin[1026] = mb1_FB1_TA1_CLKIO_N_4_mb1_FB2_BB0_CLKIO_N_2;
  assign rx_pin[1027] = mb1_FB1_TA1_CLKIO_N_5_mb1_FB2_BB0_IO_010;
  assign rx_pin[1028] = mb1_FB1_TA1_CLKIO_N_6_mb1_FB2_BB0_CLKIO_N_1;
  assign rx_pin[1029] = mb1_FB1_TA1_CLKIO_N_7_mb1_FB2_BB0_CLKIO_N_0;
  assign rx_pin[1030] = mb1_FB1_TA1_CLKIO_P_0_mb1_FB2_BB0_CLKIO_P_7;
  assign rx_pin[1031] = mb1_FB1_TA1_CLKIO_P_1_mb1_FB2_BB0_CLKIO_P_6;
  assign rx_pin[1032] = mb1_FB1_TA1_CLKIO_P_2_mb1_FB2_BB0_CLKIO_P_4;
  assign rx_pin[1033] = mb1_FB1_TA1_CLKIO_P_3_mb1_FB2_BB0_CLKIO_P_3;
  assign rx_pin[1034] = mb1_FB1_TA1_CLKIO_P_4_mb1_FB2_BB0_CLKIO_P_2;
  assign rx_pin[1035] = mb1_FB1_TA1_CLKIO_P_5_mb1_FB2_BB0_IO_011;
  assign rx_pin[1036] = mb1_FB1_TA1_CLKIO_P_6_mb1_FB2_BB0_CLKIO_P_1;
  assign rx_pin[1037] = mb1_FB1_TA1_CLKIO_P_7_mb1_FB2_BB0_CLKIO_P_0;
  assign rx_pin[1038] = mb1_FB1_TA1_IO_004_mb1_FB2_BB0_IO_006;
  assign rx_pin[1039] = mb1_FB1_TA1_IO_005_mb1_FB2_BB0_IO_007;
  assign rx_pin[1040] = mb1_FB1_TA1_IO_006_mb1_FB2_BB0_IO_004;
  assign rx_pin[1041] = mb1_FB1_TA1_IO_007_mb1_FB2_BB0_IO_005;
  assign rx_pin[1042] = mb1_FB1_TA1_IO_008_mb1_FB2_BB0_IO_022;
  assign rx_pin[1043] = mb1_FB1_TA1_IO_009_mb1_FB2_BB0_IO_023;
  assign rx_pin[1044] = mb1_FB1_TA1_IO_010_mb1_FB2_BB0_CLKIO_N_5;
  assign rx_pin[1045] = mb1_FB1_TA1_IO_011_mb1_FB2_BB0_CLKIO_P_5;
  assign rx_pin[1046] = mb1_FB1_TA1_IO_012_mb1_FB2_BB0_IO_012;
  assign rx_pin[1047] = mb1_FB1_TA1_IO_013_mb1_FB2_BB0_IO_013;
  assign rx_pin[1048] = mb1_FB1_TA1_IO_014_mb1_FB2_BB0_IO_016;
  assign rx_pin[1049] = mb1_FB1_TA1_IO_015_mb1_FB2_BB0_IO_017;
  assign rx_pin[1050] = mb1_FB1_TA1_IO_016_mb1_FB2_BB0_IO_014;
  assign rx_pin[1051] = mb1_FB1_TA1_IO_017_mb1_FB2_BB0_IO_015;
  assign rx_pin[1052] = mb1_FB1_TA1_IO_018_mb1_FB2_BB0_IO_032;
  assign rx_pin[1053] = mb1_FB1_TA1_IO_019_mb1_FB2_BB0_IO_033;
  assign rx_pin[1054] = mb1_FB1_TA1_IO_020_mb1_FB2_BB0_IO_030;
  assign rx_pin[1055] = mb1_FB1_TA1_IO_021_mb1_FB2_BB0_IO_031;
  assign rx_pin[1056] = mb1_FB1_TA1_IO_022_mb1_FB2_BB0_IO_008;
  assign rx_pin[1057] = mb1_FB1_TA1_IO_023_mb1_FB2_BB0_IO_009;
  assign rx_pin[1058] = mb1_FB1_TA1_IO_024_mb1_FB2_BB0_IO_026;
  assign rx_pin[1059] = mb1_FB1_TA1_IO_025_mb1_FB2_BB0_IO_027;
  assign rx_pin[1060] = mb1_FB1_TA1_IO_026_mb1_FB2_BB0_IO_024;
  assign rx_pin[1061] = mb1_FB1_TA1_IO_027_mb1_FB2_BB0_IO_025;
  assign rx_pin[1062] = mb1_FB1_TA1_IO_028_mb1_FB2_BB0_IO_042;
  assign rx_pin[1063] = mb1_FB1_TA1_IO_029_mb1_FB2_BB0_IO_043;
  assign rx_pin[1064] = mb1_FB1_TA1_IO_030_mb1_FB2_BB0_IO_020;
  assign rx_pin[1065] = mb1_FB1_TA1_IO_031_mb1_FB2_BB0_IO_021;
  assign rx_pin[1066] = mb1_FB1_TA1_IO_032_mb1_FB2_BB0_IO_018;
  assign rx_pin[1067] = mb1_FB1_TA1_IO_033_mb1_FB2_BB0_IO_019;
  assign rx_pin[1068] = mb1_FB1_TA1_IO_034_mb1_FB2_BB0_IO_036;
  assign rx_pin[1069] = mb1_FB1_TA1_IO_035_mb1_FB2_BB0_IO_037;
  assign rx_pin[1070] = mb1_FB1_TA1_IO_036_mb1_FB2_BB0_IO_034;
  assign rx_pin[1071] = mb1_FB1_TA1_IO_037_mb1_FB2_BB0_IO_035;
  assign rx_pin[1072] = mb1_FB1_TA1_IO_038_mb1_FB2_BB0_IO_052;
  assign rx_pin[1073] = mb1_FB1_TA1_IO_039_mb1_FB2_BB0_IO_053;
  assign rx_pin[1074] = mb1_FB1_TA1_IO_040_mb1_FB2_BB0_IO_050;
  assign rx_pin[1075] = mb1_FB1_TA1_IO_041_mb1_FB2_BB0_IO_051;
  assign rx_pin[1076] = mb1_FB1_TA1_IO_042_mb1_FB2_BB0_IO_028;
  assign rx_pin[1077] = mb1_FB1_TA1_IO_043_mb1_FB2_BB0_IO_029;
  assign rx_pin[1078] = mb1_FB1_TA1_IO_044_mb1_FB2_BB0_IO_046;
  assign rx_pin[1079] = mb1_FB1_TA1_IO_045_mb1_FB2_BB0_IO_047;
  assign rx_pin[1080] = mb1_FB1_TA1_IO_046_mb1_FB2_BB0_IO_044;
  assign rx_pin[1081] = mb1_FB1_TA1_IO_047_mb1_FB2_BB0_IO_045;
  assign rx_pin[1082] = mb1_FB1_TA1_IO_048_mb1_FB2_BB0_IO_062;
  assign rx_pin[1083] = mb1_FB1_TA1_IO_049_mb1_FB2_BB0_IO_063;
  assign rx_pin[1084] = mb1_FB1_TA1_IO_050_mb1_FB2_BB0_IO_040;
  assign rx_pin[1085] = mb1_FB1_TA1_IO_051_mb1_FB2_BB0_IO_041;
  assign rx_pin[1086] = mb1_FB1_TA1_IO_052_mb1_FB2_BB0_IO_038;
  assign rx_pin[1087] = mb1_FB1_TA1_IO_053_mb1_FB2_BB0_IO_039;
  assign rx_pin[1088] = mb1_FB1_TA1_IO_054_mb1_FB2_BB0_IO_056;
  assign rx_pin[1089] = mb1_FB1_TA1_IO_055_mb1_FB2_BB0_IO_057;
  assign rx_pin[1090] = mb1_FB1_TA1_IO_056_mb1_FB2_BB0_IO_054;
  assign rx_pin[1091] = mb1_FB1_TA1_IO_057_mb1_FB2_BB0_IO_055;
  assign rx_pin[1092] = mb1_FB1_TA1_IO_058_mb1_FB2_BB0_IO_072;
  assign rx_pin[1093] = mb1_FB1_TA1_IO_059_mb1_FB2_BB0_IO_073;
  assign rx_pin[1094] = mb1_FB1_TA1_IO_060_mb1_FB2_BB0_IO_070;
  assign rx_pin[1095] = mb1_FB1_TA1_IO_061_mb1_FB2_BB0_IO_071;
  assign rx_pin[1096] = mb1_FB1_TA1_IO_062_mb1_FB2_BB0_IO_048;
  assign rx_pin[1097] = mb1_FB1_TA1_IO_063_mb1_FB2_BB0_IO_049;
  assign rx_pin[1098] = mb1_FB1_TA1_IO_064_mb1_FB2_BB0_IO_066;
  assign rx_pin[1099] = mb1_FB1_TA1_IO_065_mb1_FB2_BB0_IO_067;
  assign rx_pin[1100] = mb1_FB1_TA1_IO_066_mb1_FB2_BB0_IO_064;
  assign rx_pin[1101] = mb1_FB1_TA1_IO_067_mb1_FB2_BB0_IO_065;
  assign rx_pin[1102] = mb1_FB1_TA1_IO_068_mb1_FB2_BB0_IO_082;
  assign rx_pin[1103] = mb1_FB1_TA1_IO_069_mb1_FB2_BB0_IO_083;
  assign rx_pin[1104] = mb1_FB1_TA1_IO_070_mb1_FB2_BB0_IO_060;
  assign rx_pin[1105] = mb1_FB1_TA1_IO_071_mb1_FB2_BB0_IO_061;
  assign rx_pin[1106] = mb1_FB1_TA1_IO_072_mb1_FB2_BB0_IO_058;
  assign rx_pin[1107] = mb1_FB1_TA1_IO_073_mb1_FB2_BB0_IO_059;
  assign rx_pin[1108] = mb1_FB1_TA1_IO_074_mb1_FB2_BB0_IO_076;
  assign rx_pin[1109] = mb1_FB1_TA1_IO_075_mb1_FB2_BB0_IO_077;
  assign rx_pin[1110] = mb1_FB1_TA1_IO_076_mb1_FB2_BB0_IO_074;
  assign rx_pin[1111] = mb1_FB1_TA1_IO_077_mb1_FB2_BB0_IO_075;
  assign rx_pin[1112] = mb1_FB1_TA1_IO_078_mb1_FB2_BB0_IO_092;
  assign rx_pin[1113] = mb1_FB1_TA1_IO_079_mb1_FB2_BB0_IO_093;
  assign rx_pin[1114] = mb1_FB1_TA1_IO_080_mb1_FB2_BB0_IO_090;
  assign rx_pin[1115] = mb1_FB1_TA1_IO_081_mb1_FB2_BB0_IO_091;
  assign rx_pin[1116] = mb1_FB1_TA1_IO_082_mb1_FB2_BB0_IO_068;
  assign rx_pin[1117] = mb1_FB1_TA1_IO_083_mb1_FB2_BB0_IO_069;
  assign rx_pin[1118] = mb1_FB1_TA1_IO_084_mb1_FB2_BB0_IO_086;
  assign rx_pin[1119] = mb1_FB1_TA1_IO_085_mb1_FB2_BB0_IO_087;
  assign rx_pin[1120] = mb1_FB1_TA1_IO_086_mb1_FB2_BB0_IO_084;
  assign rx_pin[1121] = mb1_FB1_TA1_IO_087_mb1_FB2_BB0_IO_085;
  assign rx_pin[1122] = mb1_FB1_TA1_IO_088_mb1_FB2_BB0_IO_102;
  assign rx_pin[1123] = mb1_FB1_TA1_IO_089_mb1_FB2_BB0_IO_103;
  assign rx_pin[1124] = mb1_FB1_TA1_IO_090_mb1_FB2_BB0_IO_080;
  assign rx_pin[1125] = mb1_FB1_TA1_IO_091_mb1_FB2_BB0_IO_081;
  assign rx_pin[1126] = mb1_FB1_TA1_IO_092_mb1_FB2_BB0_IO_078;
  assign rx_pin[1127] = mb1_FB1_TA1_IO_093_mb1_FB2_BB0_IO_079;
  assign rx_pin[1128] = mb1_FB1_TA1_IO_094_mb1_FB2_BB0_IO_096;
  assign rx_pin[1129] = mb1_FB1_TA1_IO_095_mb1_FB2_BB0_IO_097;
  assign rx_pin[1130] = mb1_FB1_TA1_IO_096_mb1_FB2_BB0_IO_094;
  assign rx_pin[1131] = mb1_FB1_TA1_IO_097_mb1_FB2_BB0_IO_095;
  assign rx_pin[1132] = mb1_FB1_TA1_IO_098_mb1_FB2_BB0_IO_112;
  assign rx_pin[1133] = mb1_FB1_TA1_IO_099_mb1_FB2_BB0_IO_113;
  assign rx_pin[1134] = mb1_FB1_TA1_IO_100_mb1_FB2_BB0_IO_110;
  assign rx_pin[1135] = mb1_FB1_TA1_IO_101_mb1_FB2_BB0_IO_111;
  assign rx_pin[1136] = mb1_FB1_TA1_IO_102_mb1_FB2_BB0_IO_088;
  assign rx_pin[1137] = mb1_FB1_TA1_IO_103_mb1_FB2_BB0_IO_089;
  assign rx_pin[1138] = mb1_FB1_TA1_IO_104_mb1_FB2_BB0_IO_106;
  assign rx_pin[1139] = mb1_FB1_TA1_IO_105_mb1_FB2_BB0_IO_107;
  assign rx_pin[1140] = mb1_FB1_TA1_IO_106_mb1_FB2_BB0_IO_104;
  assign rx_pin[1141] = mb1_FB1_TA1_IO_107_mb1_FB2_BB0_IO_105;
  assign rx_pin[1142] = mb1_FB1_TA1_IO_108_mb1_FB2_BB0_IO_122;
  assign rx_pin[1143] = mb1_FB1_TA1_IO_109_mb1_FB2_BB0_IO_123;
  assign rx_pin[1144] = mb1_FB1_TA1_IO_110_mb1_FB2_BB0_IO_100;
  assign rx_pin[1145] = mb1_FB1_TA1_IO_111_mb1_FB2_BB0_IO_101;
  assign rx_pin[1146] = mb1_FB1_TA1_IO_112_mb1_FB2_BB0_IO_098;
  assign rx_pin[1147] = mb1_FB1_TA1_IO_113_mb1_FB2_BB0_IO_099;
  assign rx_pin[1148] = mb1_FB1_TA1_IO_114_mb1_FB2_BB0_IO_116;
  assign rx_pin[1149] = mb1_FB1_TA1_IO_115_mb1_FB2_BB0_IO_117;
  assign rx_pin[1150] = mb1_FB1_TA1_IO_116_mb1_FB2_BB0_IO_114;
  assign rx_pin[1151] = mb1_FB1_TA1_IO_117_mb1_FB2_BB0_IO_115;
  assign rx_pin[1152] = mb1_FB1_TA1_IO_118_mb1_FB2_BB0_IO_132;
  assign rx_pin[1153] = mb1_FB1_TA1_IO_119_mb1_FB2_BB0_IO_133;
  assign rx_pin[1154] = mb1_FB1_TA1_IO_120_mb1_FB2_BB0_IO_130;
  assign rx_pin[1155] = mb1_FB1_TA1_IO_121_mb1_FB2_BB0_IO_131;
  assign rx_pin[1156] = mb1_FB1_TA1_IO_122_mb1_FB2_BB0_IO_108;
  assign rx_pin[1157] = mb1_FB1_TA1_IO_123_mb1_FB2_BB0_IO_109;
  assign rx_pin[1158] = mb1_FB1_TA1_IO_124_mb1_FB2_BB0_IO_126;
  assign rx_pin[1159] = mb1_FB1_TA1_IO_125_mb1_FB2_BB0_IO_127;
  assign rx_pin[1160] = mb1_FB1_TA1_IO_126_mb1_FB2_BB0_IO_124;
  assign rx_pin[1161] = mb1_FB1_TA1_IO_127_mb1_FB2_BB0_IO_125;
  assign rx_pin[1162] = mb1_FB1_TA1_IO_130_mb1_FB2_BB0_IO_120;
  assign rx_pin[1163] = mb1_FB1_TA1_IO_131_mb1_FB2_BB0_IO_121;
  assign rx_pin[1164] = mb1_FB1_TA1_IO_132_mb1_FB2_BB0_IO_118;
  assign rx_pin[1165] = mb1_FB1_TA1_IO_133_mb1_FB2_BB0_IO_119;
  assign rx_pin[1166] = mb1_FB1_TA1_IO_134_mb1_FB2_BB0_IO_136;
  assign rx_pin[1167] = mb1_FB1_TA1_IO_136_mb1_FB2_BB0_IO_134;
  assign rx_pin[1168] = mb1_FA1_TB2_CLKIO_N_0_mb1_FB2_BB1_CLKIO_N_7;
  assign rx_pin[1169] = mb1_FA1_TB2_CLKIO_N_1_mb1_FB2_BB1_CLKIO_N_6;
  assign rx_pin[1170] = mb1_FA1_TB2_CLKIO_N_2_mb1_FB2_BB1_CLKIO_N_4;
  assign rx_pin[1171] = mb1_FA1_TB2_CLKIO_N_3_mb1_FB2_BB1_CLKIO_N_3;
  assign rx_pin[1172] = mb1_FA1_TB2_CLKIO_N_4_mb1_FB2_BB1_CLKIO_N_2;
  assign rx_pin[1173] = mb1_FA1_TB2_CLKIO_N_5_mb1_FB2_BB1_IO_010;
  assign rx_pin[1174] = mb1_FA1_TB2_CLKIO_N_6_mb1_FB2_BB1_CLKIO_N_1;
  assign rx_pin[1175] = mb1_FA1_TB2_CLKIO_N_7_mb1_FB2_BB1_CLKIO_N_0;
  assign rx_pin[1176] = mb1_FA1_TB2_CLKIO_P_0_mb1_FB2_BB1_CLKIO_P_7;
  assign rx_pin[1177] = mb1_FA1_TB2_CLKIO_P_1_mb1_FB2_BB1_CLKIO_P_6;
  assign rx_pin[1178] = mb1_FA1_TB2_CLKIO_P_2_mb1_FB2_BB1_CLKIO_P_4;
  assign rx_pin[1179] = mb1_FA1_TB2_CLKIO_P_3_mb1_FB2_BB1_CLKIO_P_3;
  assign rx_pin[1180] = mb1_FA1_TB2_CLKIO_P_4_mb1_FB2_BB1_CLKIO_P_2;
  assign rx_pin[1181] = mb1_FA1_TB2_CLKIO_P_5_mb1_FB2_BB1_IO_011;
  assign rx_pin[1182] = mb1_FA1_TB2_CLKIO_P_6_mb1_FB2_BB1_CLKIO_P_1;
  assign rx_pin[1183] = mb1_FA1_TB2_CLKIO_P_7_mb1_FB2_BB1_CLKIO_P_0;
  assign rx_pin[1184] = mb1_FA1_TB2_IO_004_mb1_FB2_BB1_IO_006;
  assign rx_pin[1185] = mb1_FA1_TB2_IO_005_mb1_FB2_BB1_IO_007;
  assign rx_pin[1186] = mb1_FA1_TB2_IO_006_mb1_FB2_BB1_IO_004;
  assign rx_pin[1187] = mb1_FA1_TB2_IO_007_mb1_FB2_BB1_IO_005;
  assign rx_pin[1188] = mb1_FA1_TB2_IO_008_mb1_FB2_BB1_IO_022;
  assign rx_pin[1189] = mb1_FA1_TB2_IO_009_mb1_FB2_BB1_IO_023;
  assign rx_pin[1190] = mb1_FA1_TB2_IO_010_mb1_FB2_BB1_CLKIO_N_5;
  assign rx_pin[1191] = mb1_FA1_TB2_IO_011_mb1_FB2_BB1_CLKIO_P_5;
  assign rx_pin[1192] = mb1_FA1_TB2_IO_012_mb1_FB2_BB1_IO_012;
  assign rx_pin[1193] = mb1_FA1_TB2_IO_013_mb1_FB2_BB1_IO_013;
  assign rx_pin[1194] = mb1_FA1_TB2_IO_014_mb1_FB2_BB1_IO_016;
  assign rx_pin[1195] = mb1_FA1_TB2_IO_015_mb1_FB2_BB1_IO_017;
  assign rx_pin[1196] = mb1_FA1_TB2_IO_016_mb1_FB2_BB1_IO_014;
  assign rx_pin[1197] = mb1_FA1_TB2_IO_017_mb1_FB2_BB1_IO_015;
  assign rx_pin[1198] = mb1_FA1_TB2_IO_018_mb1_FB2_BB1_IO_032;
  assign rx_pin[1199] = mb1_FA1_TB2_IO_019_mb1_FB2_BB1_IO_033;
  assign rx_pin[1200] = mb1_FA1_TB2_IO_020_mb1_FB2_BB1_IO_030;
  assign rx_pin[1201] = mb1_FA1_TB2_IO_021_mb1_FB2_BB1_IO_031;
  assign rx_pin[1202] = mb1_FA1_TB2_IO_022_mb1_FB2_BB1_IO_008;
  assign rx_pin[1203] = mb1_FA1_TB2_IO_023_mb1_FB2_BB1_IO_009;
  assign rx_pin[1204] = mb1_FA1_TB2_IO_024_mb1_FB2_BB1_IO_026;
  assign rx_pin[1205] = mb1_FA1_TB2_IO_025_mb1_FB2_BB1_IO_027;
  assign rx_pin[1206] = mb1_FA1_TB2_IO_026_mb1_FB2_BB1_IO_024;
  assign rx_pin[1207] = mb1_FA1_TB2_IO_027_mb1_FB2_BB1_IO_025;
  assign rx_pin[1208] = mb1_FA1_TB2_IO_028_mb1_FB2_BB1_IO_042;
  assign rx_pin[1209] = mb1_FA1_TB2_IO_029_mb1_FB2_BB1_IO_043;
  assign rx_pin[1210] = mb1_FA1_TB2_IO_030_mb1_FB2_BB1_IO_020;
  assign rx_pin[1211] = mb1_FA1_TB2_IO_031_mb1_FB2_BB1_IO_021;
  assign rx_pin[1212] = mb1_FA1_TB2_IO_032_mb1_FB2_BB1_IO_018;
  assign rx_pin[1213] = mb1_FA1_TB2_IO_033_mb1_FB2_BB1_IO_019;
  assign rx_pin[1214] = mb1_FA1_TB2_IO_034_mb1_FB2_BB1_IO_036;
  assign rx_pin[1215] = mb1_FA1_TB2_IO_035_mb1_FB2_BB1_IO_037;
  assign rx_pin[1216] = mb1_FA1_TB2_IO_036_mb1_FB2_BB1_IO_034;
  assign rx_pin[1217] = mb1_FA1_TB2_IO_037_mb1_FB2_BB1_IO_035;
  assign rx_pin[1218] = mb1_FA1_TB2_IO_038_mb1_FB2_BB1_IO_052;
  assign rx_pin[1219] = mb1_FA1_TB2_IO_039_mb1_FB2_BB1_IO_053;
  assign rx_pin[1220] = mb1_FA1_TB2_IO_040_mb1_FB2_BB1_IO_050;
  assign rx_pin[1221] = mb1_FA1_TB2_IO_041_mb1_FB2_BB1_IO_051;
  assign rx_pin[1222] = mb1_FA1_TB2_IO_042_mb1_FB2_BB1_IO_028;
  assign rx_pin[1223] = mb1_FA1_TB2_IO_043_mb1_FB2_BB1_IO_029;
  assign rx_pin[1224] = mb1_FA1_TB2_IO_044_mb1_FB2_BB1_IO_046;
  assign rx_pin[1225] = mb1_FA1_TB2_IO_045_mb1_FB2_BB1_IO_047;
  assign rx_pin[1226] = mb1_FA1_TB2_IO_046_mb1_FB2_BB1_IO_044;
  assign rx_pin[1227] = mb1_FA1_TB2_IO_047_mb1_FB2_BB1_IO_045;
  assign rx_pin[1228] = mb1_FA1_TB2_IO_048_mb1_FB2_BB1_IO_062;
  assign rx_pin[1229] = mb1_FA1_TB2_IO_049_mb1_FB2_BB1_IO_063;
  assign rx_pin[1230] = mb1_FA1_TB2_IO_050_mb1_FB2_BB1_IO_040;
  assign rx_pin[1231] = mb1_FA1_TB2_IO_051_mb1_FB2_BB1_IO_041;
  assign rx_pin[1232] = mb1_FA1_TB2_IO_052_mb1_FB2_BB1_IO_038;
  assign rx_pin[1233] = mb1_FA1_TB2_IO_053_mb1_FB2_BB1_IO_039;
  assign rx_pin[1234] = mb1_FA1_TB2_IO_054_mb1_FB2_BB1_IO_056;
  assign rx_pin[1235] = mb1_FA1_TB2_IO_055_mb1_FB2_BB1_IO_057;
  assign rx_pin[1236] = mb1_FA1_TB2_IO_056_mb1_FB2_BB1_IO_054;
  assign rx_pin[1237] = mb1_FA1_TB2_IO_057_mb1_FB2_BB1_IO_055;
  assign rx_pin[1238] = mb1_FA1_TB2_IO_058_mb1_FB2_BB1_IO_072;
  assign rx_pin[1239] = mb1_FA1_TB2_IO_059_mb1_FB2_BB1_IO_073;
  assign rx_pin[1240] = mb1_FA1_TB2_IO_060_mb1_FB2_BB1_IO_070;
  assign rx_pin[1241] = mb1_FA1_TB2_IO_061_mb1_FB2_BB1_IO_071;
  assign rx_pin[1242] = mb1_FA1_TB2_IO_062_mb1_FB2_BB1_IO_048;
  assign rx_pin[1243] = mb1_FA1_TB2_IO_063_mb1_FB2_BB1_IO_049;
  assign rx_pin[1244] = mb1_FA1_TB2_IO_064_mb1_FB2_BB1_IO_066;
  assign rx_pin[1245] = mb1_FA1_TB2_IO_065_mb1_FB2_BB1_IO_067;
  assign rx_pin[1246] = mb1_FA1_TB2_IO_066_mb1_FB2_BB1_IO_064;
  assign rx_pin[1247] = mb1_FA1_TB2_IO_067_mb1_FB2_BB1_IO_065;
  assign rx_pin[1248] = mb1_FA1_TB2_IO_068_mb1_FB2_BB1_IO_082;
  assign rx_pin[1249] = mb1_FA1_TB2_IO_069_mb1_FB2_BB1_IO_083;
  assign rx_pin[1250] = mb1_FA1_TB2_IO_070_mb1_FB2_BB1_IO_060;
  assign rx_pin[1251] = mb1_FA1_TB2_IO_071_mb1_FB2_BB1_IO_061;
  assign rx_pin[1252] = mb1_FA1_TB2_IO_072_mb1_FB2_BB1_IO_058;
  assign rx_pin[1253] = mb1_FA1_TB2_IO_073_mb1_FB2_BB1_IO_059;
  assign rx_pin[1254] = mb1_FA1_TB2_IO_074_mb1_FB2_BB1_IO_076;
  assign rx_pin[1255] = mb1_FA1_TB2_IO_075_mb1_FB2_BB1_IO_077;
  assign rx_pin[1256] = mb1_FA1_TB2_IO_076_mb1_FB2_BB1_IO_074;
  assign rx_pin[1257] = mb1_FA1_TB2_IO_077_mb1_FB2_BB1_IO_075;
  assign rx_pin[1258] = mb1_FA1_TB2_IO_078_mb1_FB2_BB1_IO_092;
  assign rx_pin[1259] = mb1_FA1_TB2_IO_079_mb1_FB2_BB1_IO_093;
  assign rx_pin[1260] = mb1_FA1_TB2_IO_080_mb1_FB2_BB1_IO_090;
  assign rx_pin[1261] = mb1_FA1_TB2_IO_081_mb1_FB2_BB1_IO_091;
  assign rx_pin[1262] = mb1_FA1_TB2_IO_082_mb1_FB2_BB1_IO_068;
  assign rx_pin[1263] = mb1_FA1_TB2_IO_083_mb1_FB2_BB1_IO_069;
  assign rx_pin[1264] = mb1_FA1_TB2_IO_084_mb1_FB2_BB1_IO_086;
  assign rx_pin[1265] = mb1_FA1_TB2_IO_085_mb1_FB2_BB1_IO_087;
  assign rx_pin[1266] = mb1_FA1_TB2_IO_086_mb1_FB2_BB1_IO_084;
  assign rx_pin[1267] = mb1_FA1_TB2_IO_087_mb1_FB2_BB1_IO_085;
  assign rx_pin[1268] = mb1_FA1_TB2_IO_088_mb1_FB2_BB1_IO_102;
  assign rx_pin[1269] = mb1_FA1_TB2_IO_089_mb1_FB2_BB1_IO_103;
  assign rx_pin[1270] = mb1_FA1_TB2_IO_090_mb1_FB2_BB1_IO_080;
  assign rx_pin[1271] = mb1_FA1_TB2_IO_091_mb1_FB2_BB1_IO_081;
  assign rx_pin[1272] = mb1_FA1_TB2_IO_092_mb1_FB2_BB1_IO_078;
  assign rx_pin[1273] = mb1_FA1_TB2_IO_093_mb1_FB2_BB1_IO_079;
  assign rx_pin[1274] = mb1_FA1_TB2_IO_094_mb1_FB2_BB1_IO_096;
  assign rx_pin[1275] = mb1_FA1_TB2_IO_095_mb1_FB2_BB1_IO_097;
  assign rx_pin[1276] = mb1_FA1_TB2_IO_096_mb1_FB2_BB1_IO_094;
  assign rx_pin[1277] = mb1_FA1_TB2_IO_097_mb1_FB2_BB1_IO_095;
  assign rx_pin[1278] = mb1_FA1_TB2_IO_098_mb1_FB2_BB1_IO_112;
  assign rx_pin[1279] = mb1_FA1_TB2_IO_099_mb1_FB2_BB1_IO_113;
  assign rx_pin[1280] = mb1_FA1_TB2_IO_100_mb1_FB2_BB1_IO_110;
  assign rx_pin[1281] = mb1_FA1_TB2_IO_101_mb1_FB2_BB1_IO_111;
  assign rx_pin[1282] = mb1_FA1_TB2_IO_102_mb1_FB2_BB1_IO_088;
  assign rx_pin[1283] = mb1_FA1_TB2_IO_103_mb1_FB2_BB1_IO_089;
  assign rx_pin[1284] = mb1_FA1_TB2_IO_104_mb1_FB2_BB1_IO_106;
  assign rx_pin[1285] = mb1_FA1_TB2_IO_105_mb1_FB2_BB1_IO_107;
  assign rx_pin[1286] = mb1_FA1_TB2_IO_106_mb1_FB2_BB1_IO_104;
  assign rx_pin[1287] = mb1_FA1_TB2_IO_107_mb1_FB2_BB1_IO_105;
  assign rx_pin[1288] = mb1_FA1_TB2_IO_108_mb1_FB2_BB1_IO_122;
  assign rx_pin[1289] = mb1_FA1_TB2_IO_109_mb1_FB2_BB1_IO_123;
  assign rx_pin[1290] = mb1_FA1_TB2_IO_110_mb1_FB2_BB1_IO_100;
  assign rx_pin[1291] = mb1_FA1_TB2_IO_111_mb1_FB2_BB1_IO_101;
  assign rx_pin[1292] = mb1_FA1_TB2_IO_112_mb1_FB2_BB1_IO_098;
  assign rx_pin[1293] = mb1_FA1_TB2_IO_113_mb1_FB2_BB1_IO_099;
  assign rx_pin[1294] = mb1_FA1_TB2_IO_114_mb1_FB2_BB1_IO_116;
  assign rx_pin[1295] = mb1_FA1_TB2_IO_115_mb1_FB2_BB1_IO_117;
  assign rx_pin[1296] = mb1_FA1_TB2_IO_116_mb1_FB2_BB1_IO_114;
  assign rx_pin[1297] = mb1_FA1_TB2_IO_117_mb1_FB2_BB1_IO_115;
  assign rx_pin[1298] = mb1_FA1_TB2_IO_118_mb1_FB2_BB1_IO_132;
  assign rx_pin[1299] = mb1_FA1_TB2_IO_119_mb1_FB2_BB1_IO_133;
  assign rx_pin[1300] = mb1_FA1_TB2_IO_120_mb1_FB2_BB1_IO_130;
  assign rx_pin[1301] = mb1_FA1_TB2_IO_121_mb1_FB2_BB1_IO_131;
  assign rx_pin[1302] = mb1_FA1_TB2_IO_122_mb1_FB2_BB1_IO_108;
  assign rx_pin[1303] = mb1_FA1_TB2_IO_123_mb1_FB2_BB1_IO_109;
  assign rx_pin[1304] = mb1_FA1_TB2_IO_124_mb1_FB2_BB1_IO_126;
  assign rx_pin[1305] = mb1_FA1_TB2_IO_125_mb1_FB2_BB1_IO_127;
  assign rx_pin[1306] = mb1_FA1_TB2_IO_126_mb1_FB2_BB1_IO_124;
  assign rx_pin[1307] = mb1_FA1_TB2_IO_127_mb1_FB2_BB1_IO_125;
  assign rx_pin[1308] = mb1_FA1_TB2_IO_130_mb1_FB2_BB1_IO_120;
  assign rx_pin[1309] = mb1_FA1_TB2_IO_131_mb1_FB2_BB1_IO_121;
  assign rx_pin[1310] = mb1_FA1_TB2_IO_132_mb1_FB2_BB1_IO_118;
  assign rx_pin[1311] = mb1_FA1_TB2_IO_133_mb1_FB2_BB1_IO_119;
  assign rx_pin[1312] = mb1_FA1_TB2_IO_134_mb1_FB2_BB1_IO_136;
  assign rx_pin[1313] = mb1_FA1_TB2_IO_136_mb1_FB2_BB1_IO_134;
  assign rx_pin[1314] = mb1_FB1_TB0_CLKIO_N_0_mb1_FB2_BB2_CLKIO_N_7;
  assign rx_pin[1315] = mb1_FB1_TB0_CLKIO_N_1_mb1_FB2_BB2_CLKIO_N_6;
  assign rx_pin[1316] = mb1_FB1_TB0_CLKIO_N_2_mb1_FB2_BB2_CLKIO_N_4;
  assign rx_pin[1317] = mb1_FB1_TB0_CLKIO_N_3_mb1_FB2_BB2_CLKIO_N_3;
  assign rx_pin[1318] = mb1_FB1_TB0_CLKIO_N_4_mb1_FB2_BB2_CLKIO_N_2;
  assign rx_pin[1319] = mb1_FB1_TB0_CLKIO_N_5_mb1_FB2_BB2_IO_010;
  assign rx_pin[1320] = mb1_FB1_TB0_CLKIO_N_6_mb1_FB2_BB2_CLKIO_N_1;
  assign rx_pin[1321] = mb1_FB1_TB0_CLKIO_N_7_mb1_FB2_BB2_CLKIO_N_0;
  assign rx_pin[1322] = mb1_FB1_TB0_CLKIO_P_0_mb1_FB2_BB2_CLKIO_P_7;
  assign rx_pin[1323] = mb1_FB1_TB0_CLKIO_P_1_mb1_FB2_BB2_CLKIO_P_6;
  assign rx_pin[1324] = mb1_FB1_TB0_CLKIO_P_2_mb1_FB2_BB2_CLKIO_P_4;
  assign rx_pin[1325] = mb1_FB1_TB0_CLKIO_P_3_mb1_FB2_BB2_CLKIO_P_3;
  assign rx_pin[1326] = mb1_FB1_TB0_CLKIO_P_4_mb1_FB2_BB2_CLKIO_P_2;
  assign rx_pin[1327] = mb1_FB1_TB0_CLKIO_P_5_mb1_FB2_BB2_IO_011;
  assign rx_pin[1328] = mb1_FB1_TB0_CLKIO_P_6_mb1_FB2_BB2_CLKIO_P_1;
  assign rx_pin[1329] = mb1_FB1_TB0_CLKIO_P_7_mb1_FB2_BB2_CLKIO_P_0;
  assign rx_pin[1330] = mb1_FB1_TB0_IO_004_mb1_FB2_BB2_IO_006;
  assign rx_pin[1331] = mb1_FB1_TB0_IO_005_mb1_FB2_BB2_IO_007;
  assign rx_pin[1332] = mb1_FB1_TB0_IO_006_mb1_FB2_BB2_IO_004;
  assign rx_pin[1333] = mb1_FB1_TB0_IO_007_mb1_FB2_BB2_IO_005;
  assign rx_pin[1334] = mb1_FB1_TB0_IO_008_mb1_FB2_BB2_IO_022;
  assign rx_pin[1335] = mb1_FB1_TB0_IO_009_mb1_FB2_BB2_IO_023;
  assign rx_pin[1336] = mb1_FB1_TB0_IO_010_mb1_FB2_BB2_CLKIO_N_5;
  assign rx_pin[1337] = mb1_FB1_TB0_IO_011_mb1_FB2_BB2_CLKIO_P_5;
  assign rx_pin[1338] = mb1_FB1_TB0_IO_012_mb1_FB2_BB2_IO_012;
  assign rx_pin[1339] = mb1_FB1_TB0_IO_013_mb1_FB2_BB2_IO_013;
  assign rx_pin[1340] = mb1_FB1_TB0_IO_014_mb1_FB2_BB2_IO_016;
  assign rx_pin[1341] = mb1_FB1_TB0_IO_015_mb1_FB2_BB2_IO_017;
  assign rx_pin[1342] = mb1_FB1_TB0_IO_016_mb1_FB2_BB2_IO_014;
  assign rx_pin[1343] = mb1_FB1_TB0_IO_017_mb1_FB2_BB2_IO_015;
  assign rx_pin[1344] = mb1_FB1_TB0_IO_018_mb1_FB2_BB2_IO_032;
  assign rx_pin[1345] = mb1_FB1_TB0_IO_019_mb1_FB2_BB2_IO_033;
  assign rx_pin[1346] = mb1_FB1_TB0_IO_020_mb1_FB2_BB2_IO_030;
  assign rx_pin[1347] = mb1_FB1_TB0_IO_021_mb1_FB2_BB2_IO_031;
  assign rx_pin[1348] = mb1_FB1_TB0_IO_022_mb1_FB2_BB2_IO_008;
  assign rx_pin[1349] = mb1_FB1_TB0_IO_023_mb1_FB2_BB2_IO_009;
  assign rx_pin[1350] = mb1_FB1_TB0_IO_024_mb1_FB2_BB2_IO_026;
  assign rx_pin[1351] = mb1_FB1_TB0_IO_025_mb1_FB2_BB2_IO_027;
  assign rx_pin[1352] = mb1_FB1_TB0_IO_026_mb1_FB2_BB2_IO_024;
  assign rx_pin[1353] = mb1_FB1_TB0_IO_027_mb1_FB2_BB2_IO_025;
  assign rx_pin[1354] = mb1_FB1_TB0_IO_028_mb1_FB2_BB2_IO_042;
  assign rx_pin[1355] = mb1_FB1_TB0_IO_029_mb1_FB2_BB2_IO_043;
  assign rx_pin[1356] = mb1_FB1_TB0_IO_030_mb1_FB2_BB2_IO_020;
  assign rx_pin[1357] = mb1_FB1_TB0_IO_031_mb1_FB2_BB2_IO_021;
  assign rx_pin[1358] = mb1_FB1_TB0_IO_032_mb1_FB2_BB2_IO_018;
  assign rx_pin[1359] = mb1_FB1_TB0_IO_033_mb1_FB2_BB2_IO_019;
  assign rx_pin[1360] = mb1_FB1_TB0_IO_034_mb1_FB2_BB2_IO_036;
  assign rx_pin[1361] = mb1_FB1_TB0_IO_035_mb1_FB2_BB2_IO_037;
  assign rx_pin[1362] = mb1_FB1_TB0_IO_036_mb1_FB2_BB2_IO_034;
  assign rx_pin[1363] = mb1_FB1_TB0_IO_037_mb1_FB2_BB2_IO_035;
  assign rx_pin[1364] = mb1_FB1_TB0_IO_038_mb1_FB2_BB2_IO_052;
  assign rx_pin[1365] = mb1_FB1_TB0_IO_039_mb1_FB2_BB2_IO_053;
  assign rx_pin[1366] = mb1_FB1_TB0_IO_040_mb1_FB2_BB2_IO_050;
  assign rx_pin[1367] = mb1_FB1_TB0_IO_041_mb1_FB2_BB2_IO_051;
  assign rx_pin[1368] = mb1_FB1_TB0_IO_042_mb1_FB2_BB2_IO_028;
  assign rx_pin[1369] = mb1_FB1_TB0_IO_043_mb1_FB2_BB2_IO_029;
  assign rx_pin[1370] = mb1_FB1_TB0_IO_044_mb1_FB2_BB2_IO_046;
  assign rx_pin[1371] = mb1_FB1_TB0_IO_045_mb1_FB2_BB2_IO_047;
  assign rx_pin[1372] = mb1_FB1_TB0_IO_046_mb1_FB2_BB2_IO_044;
  assign rx_pin[1373] = mb1_FB1_TB0_IO_047_mb1_FB2_BB2_IO_045;
  assign rx_pin[1374] = mb1_FB1_TB0_IO_048_mb1_FB2_BB2_IO_062;
  assign rx_pin[1375] = mb1_FB1_TB0_IO_049_mb1_FB2_BB2_IO_063;
  assign rx_pin[1376] = mb1_FB1_TB0_IO_050_mb1_FB2_BB2_IO_040;
  assign rx_pin[1377] = mb1_FB1_TB0_IO_051_mb1_FB2_BB2_IO_041;
  assign rx_pin[1378] = mb1_FB1_TB0_IO_052_mb1_FB2_BB2_IO_038;
  assign rx_pin[1379] = mb1_FB1_TB0_IO_053_mb1_FB2_BB2_IO_039;
  assign rx_pin[1380] = mb1_FB1_TB0_IO_054_mb1_FB2_BB2_IO_056;
  assign rx_pin[1381] = mb1_FB1_TB0_IO_055_mb1_FB2_BB2_IO_057;
  assign rx_pin[1382] = mb1_FB1_TB0_IO_056_mb1_FB2_BB2_IO_054;
  assign rx_pin[1383] = mb1_FB1_TB0_IO_057_mb1_FB2_BB2_IO_055;
  assign rx_pin[1384] = mb1_FB1_TB0_IO_058_mb1_FB2_BB2_IO_072;
  assign rx_pin[1385] = mb1_FB1_TB0_IO_059_mb1_FB2_BB2_IO_073;
  assign rx_pin[1386] = mb1_FB1_TB0_IO_060_mb1_FB2_BB2_IO_070;
  assign rx_pin[1387] = mb1_FB1_TB0_IO_061_mb1_FB2_BB2_IO_071;
  assign rx_pin[1388] = mb1_FB1_TB0_IO_062_mb1_FB2_BB2_IO_048;
  assign rx_pin[1389] = mb1_FB1_TB0_IO_063_mb1_FB2_BB2_IO_049;
  assign rx_pin[1390] = mb1_FB1_TB0_IO_064_mb1_FB2_BB2_IO_066;
  assign rx_pin[1391] = mb1_FB1_TB0_IO_065_mb1_FB2_BB2_IO_067;
  assign rx_pin[1392] = mb1_FB1_TB0_IO_066_mb1_FB2_BB2_IO_064;
  assign rx_pin[1393] = mb1_FB1_TB0_IO_067_mb1_FB2_BB2_IO_065;
  assign rx_pin[1394] = mb1_FB1_TB0_IO_068_mb1_FB2_BB2_IO_082;
  assign rx_pin[1395] = mb1_FB1_TB0_IO_069_mb1_FB2_BB2_IO_083;
  assign rx_pin[1396] = mb1_FB1_TB0_IO_070_mb1_FB2_BB2_IO_060;
  assign rx_pin[1397] = mb1_FB1_TB0_IO_071_mb1_FB2_BB2_IO_061;
  assign rx_pin[1398] = mb1_FB1_TB0_IO_072_mb1_FB2_BB2_IO_058;
  assign rx_pin[1399] = mb1_FB1_TB0_IO_073_mb1_FB2_BB2_IO_059;
  assign rx_pin[1400] = mb1_FB1_TB0_IO_074_mb1_FB2_BB2_IO_076;
  assign rx_pin[1401] = mb1_FB1_TB0_IO_075_mb1_FB2_BB2_IO_077;
  assign rx_pin[1402] = mb1_FB1_TB0_IO_076_mb1_FB2_BB2_IO_074;
  assign rx_pin[1403] = mb1_FB1_TB0_IO_077_mb1_FB2_BB2_IO_075;
  assign rx_pin[1404] = mb1_FB1_TB0_IO_078_mb1_FB2_BB2_IO_092;
  assign rx_pin[1405] = mb1_FB1_TB0_IO_079_mb1_FB2_BB2_IO_093;
  assign rx_pin[1406] = mb1_FB1_TB0_IO_080_mb1_FB2_BB2_IO_090;
  assign rx_pin[1407] = mb1_FB1_TB0_IO_081_mb1_FB2_BB2_IO_091;
  assign rx_pin[1408] = mb1_FB1_TB0_IO_082_mb1_FB2_BB2_IO_068;
  assign rx_pin[1409] = mb1_FB1_TB0_IO_083_mb1_FB2_BB2_IO_069;
  assign rx_pin[1410] = mb1_FB1_TB0_IO_084_mb1_FB2_BB2_IO_086;
  assign rx_pin[1411] = mb1_FB1_TB0_IO_085_mb1_FB2_BB2_IO_087;
  assign rx_pin[1412] = mb1_FB1_TB0_IO_086_mb1_FB2_BB2_IO_084;
  assign rx_pin[1413] = mb1_FB1_TB0_IO_087_mb1_FB2_BB2_IO_085;
  assign rx_pin[1414] = mb1_FB1_TB0_IO_088_mb1_FB2_BB2_IO_102;
  assign rx_pin[1415] = mb1_FB1_TB0_IO_089_mb1_FB2_BB2_IO_103;
  assign rx_pin[1416] = mb1_FB1_TB0_IO_090_mb1_FB2_BB2_IO_080;
  assign rx_pin[1417] = mb1_FB1_TB0_IO_091_mb1_FB2_BB2_IO_081;
  assign rx_pin[1418] = mb1_FB1_TB0_IO_092_mb1_FB2_BB2_IO_078;
  assign rx_pin[1419] = mb1_FB1_TB0_IO_093_mb1_FB2_BB2_IO_079;
  assign rx_pin[1420] = mb1_FB1_TB0_IO_094_mb1_FB2_BB2_IO_096;
  assign rx_pin[1421] = mb1_FB1_TB0_IO_095_mb1_FB2_BB2_IO_097;
  assign rx_pin[1422] = mb1_FB1_TB0_IO_096_mb1_FB2_BB2_IO_094;
  assign rx_pin[1423] = mb1_FB1_TB0_IO_097_mb1_FB2_BB2_IO_095;
  assign rx_pin[1424] = mb1_FB1_TB0_IO_098_mb1_FB2_BB2_IO_112;
  assign rx_pin[1425] = mb1_FB1_TB0_IO_099_mb1_FB2_BB2_IO_113;
  assign rx_pin[1426] = mb1_FB1_TB0_IO_100_mb1_FB2_BB2_IO_110;
  assign rx_pin[1427] = mb1_FB1_TB0_IO_101_mb1_FB2_BB2_IO_111;
  assign rx_pin[1428] = mb1_FB1_TB0_IO_102_mb1_FB2_BB2_IO_088;
  assign rx_pin[1429] = mb1_FB1_TB0_IO_103_mb1_FB2_BB2_IO_089;
  assign rx_pin[1430] = mb1_FB1_TB0_IO_104_mb1_FB2_BB2_IO_106;
  assign rx_pin[1431] = mb1_FB1_TB0_IO_105_mb1_FB2_BB2_IO_107;
  assign rx_pin[1432] = mb1_FB1_TB0_IO_106_mb1_FB2_BB2_IO_104;
  assign rx_pin[1433] = mb1_FB1_TB0_IO_107_mb1_FB2_BB2_IO_105;
  assign rx_pin[1434] = mb1_FB1_TB0_IO_108_mb1_FB2_BB2_IO_122;
  assign rx_pin[1435] = mb1_FB1_TB0_IO_109_mb1_FB2_BB2_IO_123;
  assign rx_pin[1436] = mb1_FB1_TB0_IO_110_mb1_FB2_BB2_IO_100;
  assign rx_pin[1437] = mb1_FB1_TB0_IO_111_mb1_FB2_BB2_IO_101;
  assign rx_pin[1438] = mb1_FB1_TB0_IO_112_mb1_FB2_BB2_IO_098;
  assign rx_pin[1439] = mb1_FB1_TB0_IO_113_mb1_FB2_BB2_IO_099;
  assign rx_pin[1440] = mb1_FB1_TB0_IO_114_mb1_FB2_BB2_IO_116;
  assign rx_pin[1441] = mb1_FB1_TB0_IO_115_mb1_FB2_BB2_IO_117;
  assign rx_pin[1442] = mb1_FB1_TB0_IO_116_mb1_FB2_BB2_IO_114;
  assign rx_pin[1443] = mb1_FB1_TB0_IO_117_mb1_FB2_BB2_IO_115;
  assign rx_pin[1444] = mb1_FB1_TB0_IO_118_mb1_FB2_BB2_IO_132;
  assign rx_pin[1445] = mb1_FB1_TB0_IO_119_mb1_FB2_BB2_IO_133;
  assign rx_pin[1446] = mb1_FB1_TB0_IO_120_mb1_FB2_BB2_IO_130;
  assign rx_pin[1447] = mb1_FB1_TB0_IO_121_mb1_FB2_BB2_IO_131;
  assign rx_pin[1448] = mb1_FB1_TB0_IO_122_mb1_FB2_BB2_IO_108;
  assign rx_pin[1449] = mb1_FB1_TB0_IO_123_mb1_FB2_BB2_IO_109;
  assign rx_pin[1450] = mb1_FB1_TB0_IO_124_mb1_FB2_BB2_IO_126;
  assign rx_pin[1451] = mb1_FB1_TB0_IO_125_mb1_FB2_BB2_IO_127;
  assign rx_pin[1452] = mb1_FB1_TB0_IO_126_mb1_FB2_BB2_IO_124;
  assign rx_pin[1453] = mb1_FB1_TB0_IO_127_mb1_FB2_BB2_IO_125;
  assign rx_pin[1454] = mb1_FB1_TB0_IO_130_mb1_FB2_BB2_IO_120;
  assign rx_pin[1455] = mb1_FB1_TB0_IO_131_mb1_FB2_BB2_IO_121;
  assign rx_pin[1456] = mb1_FB1_TB0_IO_132_mb1_FB2_BB2_IO_118;
  assign rx_pin[1457] = mb1_FB1_TB0_IO_133_mb1_FB2_BB2_IO_119;
  assign rx_pin[1458] = mb1_FB1_TB0_IO_134_mb1_FB2_BB2_IO_136;
  assign rx_pin[1459] = mb1_FB1_TB0_IO_136_mb1_FB2_BB2_IO_134;

  dbst # (
    .DEVICE             ( "XVUP"   ),
    .TX_PINS            ( TX_PINS               ),
    .RX_PINS            ( RX_PINS               ),
    .DIFF_ENABLED       ( 0 ),
    .USE_CLK_INPUT_BUFG ( USE_CLK_INPUT_BUFG    )
  ) U_DBST (
    .tx_pin        (             ),
    .tx_pin_p      (             ),
    .tx_pin_n      (             ),
    .rx_pin        ( rx_pin      ),
    .rx_pin_p      ( '0          ),
    .rx_pin_n      ( '0          ),
    .clk_p         ( CLK_P[1:0]  ),
    .clk_n         ( CLK_N[1:0]  ),
    .sync_p        ( SYNC_P[1:0] ),
    .sync_n        ( SYNC_N[1:0] ),
    .dmbi_f2h_o    ( DMBI_F2H    ),
    .dmbi_h2f_i    ( DMBI_H2F    )
  );
  
endmodule
