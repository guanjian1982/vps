// Unpublished work. Copyright 2022 Siemens                         
// This material contains trade secrets or otherwise                
// confidential information owned by Siemens Industry Software Inc. 
// or its affiliates (collectively, "SISW"), or its licensors.      
// Access to and use of this information is strictly limited as     
// set forth in the Customer's applicable agreements with SISW.     
// This file was generated by profpga_brdgen version 14.0 
//   on Fri Dec 15 16:10:03 2023 

`timescale 1 ps / 1 ps

// Disable implicit declaration of wires
`default_nettype none

module top_fpga_mb1fb1
   (
    input  wire [7:0]  CLK_N,
    input  wire [7:0]  CLK_P,
    input  wire [7:0]  SYNC_N,
    input  wire [7:0]  SYNC_P,
    output wire [3:0]  SRC_CLK_N,
    output wire [3:0]  SRC_CLK_P,
    output wire [3:0]  SRC_SYNC_N,
    output wire [3:0]  SRC_SYNC_P,
    output wire [19:0] DMBI_F2H,
    input  wire [19:0] DMBI_H2F,
    output wire        mb1_FB1_TA1_CLKIO_N_0_mb1_FB2_BB0_CLKIO_N_7,
    output wire        mb1_FB1_TA1_CLKIO_N_1_mb1_FB2_BB0_CLKIO_N_6,
    output wire        mb1_FB1_TA1_CLKIO_N_2_mb1_FB2_BB0_CLKIO_N_4,
    output wire        mb1_FB1_TA1_CLKIO_N_3_mb1_FB2_BB0_CLKIO_N_3,
    output wire        mb1_FB1_TA1_CLKIO_N_4_mb1_FB2_BB0_CLKIO_N_2,
    output wire        mb1_FB1_TA1_CLKIO_N_5_mb1_FB2_BB0_IO_010,
    output wire        mb1_FB1_TA1_CLKIO_N_6_mb1_FB2_BB0_CLKIO_N_1,
    output wire        mb1_FB1_TA1_CLKIO_N_7_mb1_FB2_BB0_CLKIO_N_0,
    output wire        mb1_FB1_TA1_CLKIO_P_0_mb1_FB2_BB0_CLKIO_P_7,
    output wire        mb1_FB1_TA1_CLKIO_P_1_mb1_FB2_BB0_CLKIO_P_6,
    output wire        mb1_FB1_TA1_CLKIO_P_2_mb1_FB2_BB0_CLKIO_P_4,
    output wire        mb1_FB1_TA1_CLKIO_P_3_mb1_FB2_BB0_CLKIO_P_3,
    output wire        mb1_FB1_TA1_CLKIO_P_4_mb1_FB2_BB0_CLKIO_P_2,
    output wire        mb1_FB1_TA1_CLKIO_P_5_mb1_FB2_BB0_IO_011,
    output wire        mb1_FB1_TA1_CLKIO_P_6_mb1_FB2_BB0_CLKIO_P_1,
    output wire        mb1_FB1_TA1_CLKIO_P_7_mb1_FB2_BB0_CLKIO_P_0,
    output wire        mb1_FB1_TA1_IO_004_mb1_FB2_BB0_IO_006,
    output wire        mb1_FB1_TA1_IO_005_mb1_FB2_BB0_IO_007,
    output wire        mb1_FB1_TA1_IO_006_mb1_FB2_BB0_IO_004,
    output wire        mb1_FB1_TA1_IO_007_mb1_FB2_BB0_IO_005,
    output wire        mb1_FB1_TA1_IO_008_mb1_FB2_BB0_IO_022,
    output wire        mb1_FB1_TA1_IO_009_mb1_FB2_BB0_IO_023,
    output wire        mb1_FB1_TA1_IO_010_mb1_FB2_BB0_CLKIO_N_5,
    output wire        mb1_FB1_TA1_IO_011_mb1_FB2_BB0_CLKIO_P_5,
    output wire        mb1_FB1_TA1_IO_012_mb1_FB2_BB0_IO_012,
    output wire        mb1_FB1_TA1_IO_013_mb1_FB2_BB0_IO_013,
    output wire        mb1_FB1_TA1_IO_014_mb1_FB2_BB0_IO_016,
    output wire        mb1_FB1_TA1_IO_015_mb1_FB2_BB0_IO_017,
    output wire        mb1_FB1_TA1_IO_016_mb1_FB2_BB0_IO_014,
    output wire        mb1_FB1_TA1_IO_017_mb1_FB2_BB0_IO_015,
    output wire        mb1_FB1_TA1_IO_018_mb1_FB2_BB0_IO_032,
    output wire        mb1_FB1_TA1_IO_019_mb1_FB2_BB0_IO_033,
    output wire        mb1_FB1_TA1_IO_020_mb1_FB2_BB0_IO_030,
    output wire        mb1_FB1_TA1_IO_021_mb1_FB2_BB0_IO_031,
    output wire        mb1_FB1_TA1_IO_022_mb1_FB2_BB0_IO_008,
    output wire        mb1_FB1_TA1_IO_023_mb1_FB2_BB0_IO_009,
    output wire        mb1_FB1_TA1_IO_024_mb1_FB2_BB0_IO_026,
    output wire        mb1_FB1_TA1_IO_025_mb1_FB2_BB0_IO_027,
    output wire        mb1_FB1_TA1_IO_026_mb1_FB2_BB0_IO_024,
    output wire        mb1_FB1_TA1_IO_027_mb1_FB2_BB0_IO_025,
    output wire        mb1_FB1_TA1_IO_028_mb1_FB2_BB0_IO_042,
    output wire        mb1_FB1_TA1_IO_029_mb1_FB2_BB0_IO_043,
    output wire        mb1_FB1_TA1_IO_030_mb1_FB2_BB0_IO_020,
    output wire        mb1_FB1_TA1_IO_031_mb1_FB2_BB0_IO_021,
    output wire        mb1_FB1_TA1_IO_032_mb1_FB2_BB0_IO_018,
    output wire        mb1_FB1_TA1_IO_033_mb1_FB2_BB0_IO_019,
    output wire        mb1_FB1_TA1_IO_034_mb1_FB2_BB0_IO_036,
    output wire        mb1_FB1_TA1_IO_035_mb1_FB2_BB0_IO_037,
    output wire        mb1_FB1_TA1_IO_036_mb1_FB2_BB0_IO_034,
    output wire        mb1_FB1_TA1_IO_037_mb1_FB2_BB0_IO_035,
    output wire        mb1_FB1_TA1_IO_038_mb1_FB2_BB0_IO_052,
    output wire        mb1_FB1_TA1_IO_039_mb1_FB2_BB0_IO_053,
    output wire        mb1_FB1_TA1_IO_040_mb1_FB2_BB0_IO_050,
    output wire        mb1_FB1_TA1_IO_041_mb1_FB2_BB0_IO_051,
    output wire        mb1_FB1_TA1_IO_042_mb1_FB2_BB0_IO_028,
    output wire        mb1_FB1_TA1_IO_043_mb1_FB2_BB0_IO_029,
    output wire        mb1_FB1_TA1_IO_044_mb1_FB2_BB0_IO_046,
    output wire        mb1_FB1_TA1_IO_045_mb1_FB2_BB0_IO_047,
    output wire        mb1_FB1_TA1_IO_046_mb1_FB2_BB0_IO_044,
    output wire        mb1_FB1_TA1_IO_047_mb1_FB2_BB0_IO_045,
    output wire        mb1_FB1_TA1_IO_048_mb1_FB2_BB0_IO_062,
    output wire        mb1_FB1_TA1_IO_049_mb1_FB2_BB0_IO_063,
    output wire        mb1_FB1_TA1_IO_050_mb1_FB2_BB0_IO_040,
    output wire        mb1_FB1_TA1_IO_051_mb1_FB2_BB0_IO_041,
    output wire        mb1_FB1_TA1_IO_052_mb1_FB2_BB0_IO_038,
    output wire        mb1_FB1_TA1_IO_053_mb1_FB2_BB0_IO_039,
    output wire        mb1_FB1_TA1_IO_054_mb1_FB2_BB0_IO_056,
    output wire        mb1_FB1_TA1_IO_055_mb1_FB2_BB0_IO_057,
    output wire        mb1_FB1_TA1_IO_056_mb1_FB2_BB0_IO_054,
    output wire        mb1_FB1_TA1_IO_057_mb1_FB2_BB0_IO_055,
    output wire        mb1_FB1_TA1_IO_058_mb1_FB2_BB0_IO_072,
    output wire        mb1_FB1_TA1_IO_059_mb1_FB2_BB0_IO_073,
    output wire        mb1_FB1_TA1_IO_060_mb1_FB2_BB0_IO_070,
    output wire        mb1_FB1_TA1_IO_061_mb1_FB2_BB0_IO_071,
    output wire        mb1_FB1_TA1_IO_062_mb1_FB2_BB0_IO_048,
    output wire        mb1_FB1_TA1_IO_063_mb1_FB2_BB0_IO_049,
    output wire        mb1_FB1_TA1_IO_064_mb1_FB2_BB0_IO_066,
    output wire        mb1_FB1_TA1_IO_065_mb1_FB2_BB0_IO_067,
    output wire        mb1_FB1_TA1_IO_066_mb1_FB2_BB0_IO_064,
    output wire        mb1_FB1_TA1_IO_067_mb1_FB2_BB0_IO_065,
    output wire        mb1_FB1_TA1_IO_068_mb1_FB2_BB0_IO_082,
    output wire        mb1_FB1_TA1_IO_069_mb1_FB2_BB0_IO_083,
    output wire        mb1_FB1_TA1_IO_070_mb1_FB2_BB0_IO_060,
    output wire        mb1_FB1_TA1_IO_071_mb1_FB2_BB0_IO_061,
    output wire        mb1_FB1_TA1_IO_072_mb1_FB2_BB0_IO_058,
    output wire        mb1_FB1_TA1_IO_073_mb1_FB2_BB0_IO_059,
    output wire        mb1_FB1_TA1_IO_074_mb1_FB2_BB0_IO_076,
    output wire        mb1_FB1_TA1_IO_075_mb1_FB2_BB0_IO_077,
    output wire        mb1_FB1_TA1_IO_076_mb1_FB2_BB0_IO_074,
    output wire        mb1_FB1_TA1_IO_077_mb1_FB2_BB0_IO_075,
    output wire        mb1_FB1_TA1_IO_078_mb1_FB2_BB0_IO_092,
    output wire        mb1_FB1_TA1_IO_079_mb1_FB2_BB0_IO_093,
    output wire        mb1_FB1_TA1_IO_080_mb1_FB2_BB0_IO_090,
    output wire        mb1_FB1_TA1_IO_081_mb1_FB2_BB0_IO_091,
    output wire        mb1_FB1_TA1_IO_082_mb1_FB2_BB0_IO_068,
    output wire        mb1_FB1_TA1_IO_083_mb1_FB2_BB0_IO_069,
    output wire        mb1_FB1_TA1_IO_084_mb1_FB2_BB0_IO_086,
    output wire        mb1_FB1_TA1_IO_085_mb1_FB2_BB0_IO_087,
    output wire        mb1_FB1_TA1_IO_086_mb1_FB2_BB0_IO_084,
    output wire        mb1_FB1_TA1_IO_087_mb1_FB2_BB0_IO_085,
    output wire        mb1_FB1_TA1_IO_088_mb1_FB2_BB0_IO_102,
    output wire        mb1_FB1_TA1_IO_089_mb1_FB2_BB0_IO_103,
    output wire        mb1_FB1_TA1_IO_090_mb1_FB2_BB0_IO_080,
    output wire        mb1_FB1_TA1_IO_091_mb1_FB2_BB0_IO_081,
    output wire        mb1_FB1_TA1_IO_092_mb1_FB2_BB0_IO_078,
    output wire        mb1_FB1_TA1_IO_093_mb1_FB2_BB0_IO_079,
    output wire        mb1_FB1_TA1_IO_094_mb1_FB2_BB0_IO_096,
    output wire        mb1_FB1_TA1_IO_095_mb1_FB2_BB0_IO_097,
    output wire        mb1_FB1_TA1_IO_096_mb1_FB2_BB0_IO_094,
    output wire        mb1_FB1_TA1_IO_097_mb1_FB2_BB0_IO_095,
    output wire        mb1_FB1_TA1_IO_098_mb1_FB2_BB0_IO_112,
    output wire        mb1_FB1_TA1_IO_099_mb1_FB2_BB0_IO_113,
    output wire        mb1_FB1_TA1_IO_100_mb1_FB2_BB0_IO_110,
    output wire        mb1_FB1_TA1_IO_101_mb1_FB2_BB0_IO_111,
    output wire        mb1_FB1_TA1_IO_102_mb1_FB2_BB0_IO_088,
    output wire        mb1_FB1_TA1_IO_103_mb1_FB2_BB0_IO_089,
    output wire        mb1_FB1_TA1_IO_104_mb1_FB2_BB0_IO_106,
    output wire        mb1_FB1_TA1_IO_105_mb1_FB2_BB0_IO_107,
    output wire        mb1_FB1_TA1_IO_106_mb1_FB2_BB0_IO_104,
    output wire        mb1_FB1_TA1_IO_107_mb1_FB2_BB0_IO_105,
    output wire        mb1_FB1_TA1_IO_108_mb1_FB2_BB0_IO_122,
    output wire        mb1_FB1_TA1_IO_109_mb1_FB2_BB0_IO_123,
    output wire        mb1_FB1_TA1_IO_110_mb1_FB2_BB0_IO_100,
    output wire        mb1_FB1_TA1_IO_111_mb1_FB2_BB0_IO_101,
    output wire        mb1_FB1_TA1_IO_112_mb1_FB2_BB0_IO_098,
    output wire        mb1_FB1_TA1_IO_113_mb1_FB2_BB0_IO_099,
    output wire        mb1_FB1_TA1_IO_114_mb1_FB2_BB0_IO_116,
    output wire        mb1_FB1_TA1_IO_115_mb1_FB2_BB0_IO_117,
    output wire        mb1_FB1_TA1_IO_116_mb1_FB2_BB0_IO_114,
    output wire        mb1_FB1_TA1_IO_117_mb1_FB2_BB0_IO_115,
    output wire        mb1_FB1_TA1_IO_118_mb1_FB2_BB0_IO_132,
    output wire        mb1_FB1_TA1_IO_119_mb1_FB2_BB0_IO_133,
    output wire        mb1_FB1_TA1_IO_120_mb1_FB2_BB0_IO_130,
    output wire        mb1_FB1_TA1_IO_121_mb1_FB2_BB0_IO_131,
    output wire        mb1_FB1_TA1_IO_122_mb1_FB2_BB0_IO_108,
    output wire        mb1_FB1_TA1_IO_123_mb1_FB2_BB0_IO_109,
    output wire        mb1_FB1_TA1_IO_124_mb1_FB2_BB0_IO_126,
    output wire        mb1_FB1_TA1_IO_125_mb1_FB2_BB0_IO_127,
    output wire        mb1_FB1_TA1_IO_126_mb1_FB2_BB0_IO_124,
    output wire        mb1_FB1_TA1_IO_127_mb1_FB2_BB0_IO_125,
    output wire        mb1_FB1_TA1_IO_130_mb1_FB2_BB0_IO_120,
    output wire        mb1_FB1_TA1_IO_131_mb1_FB2_BB0_IO_121,
    output wire        mb1_FB1_TA1_IO_132_mb1_FB2_BB0_IO_118,
    output wire        mb1_FB1_TA1_IO_133_mb1_FB2_BB0_IO_119,
    output wire        mb1_FB1_TA1_IO_134_mb1_FB2_BB0_IO_136,
    output wire        mb1_FB1_TA1_IO_136_mb1_FB2_BB0_IO_134,
    input wire        mb1_FA1_TA1_CLKIO_N_0_mb1_FB1_TA2_CLKIO_N_7,
    input wire        mb1_FA1_TA1_CLKIO_N_1_mb1_FB1_TA2_CLKIO_N_6,
    input wire        mb1_FA1_TA1_CLKIO_N_2_mb1_FB1_TA2_CLKIO_N_4,
    input wire        mb1_FA1_TA1_CLKIO_N_3_mb1_FB1_TA2_CLKIO_N_3,
    input wire        mb1_FA1_TA1_CLKIO_N_4_mb1_FB1_TA2_CLKIO_N_2,
    input wire        mb1_FA1_TA1_CLKIO_N_5_mb1_FB1_TA2_IO_010,
    input wire        mb1_FA1_TA1_CLKIO_N_6_mb1_FB1_TA2_CLKIO_N_1,
    input wire        mb1_FA1_TA1_CLKIO_N_7_mb1_FB1_TA2_CLKIO_N_0,
    input wire        mb1_FA1_TA1_CLKIO_P_0_mb1_FB1_TA2_CLKIO_P_7,
    input wire        mb1_FA1_TA1_CLKIO_P_1_mb1_FB1_TA2_CLKIO_P_6,
    input wire        mb1_FA1_TA1_CLKIO_P_2_mb1_FB1_TA2_CLKIO_P_4,
    input wire        mb1_FA1_TA1_CLKIO_P_3_mb1_FB1_TA2_CLKIO_P_3,
    input wire        mb1_FA1_TA1_CLKIO_P_4_mb1_FB1_TA2_CLKIO_P_2,
    input wire        mb1_FA1_TA1_CLKIO_P_5_mb1_FB1_TA2_IO_011,
    input wire        mb1_FA1_TA1_CLKIO_P_6_mb1_FB1_TA2_CLKIO_P_1,
    input wire        mb1_FA1_TA1_CLKIO_P_7_mb1_FB1_TA2_CLKIO_P_0,
    input wire        mb1_FA1_TA1_IO_004_mb1_FB1_TA2_IO_006,
    input wire        mb1_FA1_TA1_IO_005_mb1_FB1_TA2_IO_007,
    input wire        mb1_FA1_TA1_IO_006_mb1_FB1_TA2_IO_004,
    input wire        mb1_FA1_TA1_IO_007_mb1_FB1_TA2_IO_005,
    input wire        mb1_FA1_TA1_IO_008_mb1_FB1_TA2_IO_022,
    input wire        mb1_FA1_TA1_IO_009_mb1_FB1_TA2_IO_023,
    input wire        mb1_FA1_TA1_IO_010_mb1_FB1_TA2_CLKIO_N_5,
    input wire        mb1_FA1_TA1_IO_011_mb1_FB1_TA2_CLKIO_P_5,
    input wire        mb1_FA1_TA1_IO_012_mb1_FB1_TA2_IO_012,
    input wire        mb1_FA1_TA1_IO_013_mb1_FB1_TA2_IO_013,
    input wire        mb1_FA1_TA1_IO_014_mb1_FB1_TA2_IO_016,
    input wire        mb1_FA1_TA1_IO_015_mb1_FB1_TA2_IO_017,
    input wire        mb1_FA1_TA1_IO_016_mb1_FB1_TA2_IO_014,
    input wire        mb1_FA1_TA1_IO_017_mb1_FB1_TA2_IO_015,
    input wire        mb1_FA1_TA1_IO_018_mb1_FB1_TA2_IO_032,
    input wire        mb1_FA1_TA1_IO_019_mb1_FB1_TA2_IO_033,
    input wire        mb1_FA1_TA1_IO_020_mb1_FB1_TA2_IO_030,
    input wire        mb1_FA1_TA1_IO_021_mb1_FB1_TA2_IO_031,
    input wire        mb1_FA1_TA1_IO_022_mb1_FB1_TA2_IO_008,
    input wire        mb1_FA1_TA1_IO_023_mb1_FB1_TA2_IO_009,
    input wire        mb1_FA1_TA1_IO_024_mb1_FB1_TA2_IO_026,
    input wire        mb1_FA1_TA1_IO_025_mb1_FB1_TA2_IO_027,
    input wire        mb1_FA1_TA1_IO_026_mb1_FB1_TA2_IO_024,
    input wire        mb1_FA1_TA1_IO_027_mb1_FB1_TA2_IO_025,
    input wire        mb1_FA1_TA1_IO_028_mb1_FB1_TA2_IO_042,
    input wire        mb1_FA1_TA1_IO_029_mb1_FB1_TA2_IO_043,
    input wire        mb1_FA1_TA1_IO_030_mb1_FB1_TA2_IO_020,
    input wire        mb1_FA1_TA1_IO_031_mb1_FB1_TA2_IO_021,
    input wire        mb1_FA1_TA1_IO_032_mb1_FB1_TA2_IO_018,
    input wire        mb1_FA1_TA1_IO_033_mb1_FB1_TA2_IO_019,
    input wire        mb1_FA1_TA1_IO_034_mb1_FB1_TA2_IO_036,
    input wire        mb1_FA1_TA1_IO_035_mb1_FB1_TA2_IO_037,
    input wire        mb1_FA1_TA1_IO_036_mb1_FB1_TA2_IO_034,
    input wire        mb1_FA1_TA1_IO_037_mb1_FB1_TA2_IO_035,
    input wire        mb1_FA1_TA1_IO_038_mb1_FB1_TA2_IO_052,
    input wire        mb1_FA1_TA1_IO_039_mb1_FB1_TA2_IO_053,
    input wire        mb1_FA1_TA1_IO_040_mb1_FB1_TA2_IO_050,
    input wire        mb1_FA1_TA1_IO_041_mb1_FB1_TA2_IO_051,
    input wire        mb1_FA1_TA1_IO_042_mb1_FB1_TA2_IO_028,
    input wire        mb1_FA1_TA1_IO_043_mb1_FB1_TA2_IO_029,
    input wire        mb1_FA1_TA1_IO_044_mb1_FB1_TA2_IO_046,
    input wire        mb1_FA1_TA1_IO_045_mb1_FB1_TA2_IO_047,
    input wire        mb1_FA1_TA1_IO_046_mb1_FB1_TA2_IO_044,
    input wire        mb1_FA1_TA1_IO_047_mb1_FB1_TA2_IO_045,
    input wire        mb1_FA1_TA1_IO_048_mb1_FB1_TA2_IO_062,
    input wire        mb1_FA1_TA1_IO_049_mb1_FB1_TA2_IO_063,
    input wire        mb1_FA1_TA1_IO_050_mb1_FB1_TA2_IO_040,
    input wire        mb1_FA1_TA1_IO_051_mb1_FB1_TA2_IO_041,
    input wire        mb1_FA1_TA1_IO_052_mb1_FB1_TA2_IO_038,
    input wire        mb1_FA1_TA1_IO_053_mb1_FB1_TA2_IO_039,
    input wire        mb1_FA1_TA1_IO_054_mb1_FB1_TA2_IO_056,
    input wire        mb1_FA1_TA1_IO_055_mb1_FB1_TA2_IO_057,
    input wire        mb1_FA1_TA1_IO_056_mb1_FB1_TA2_IO_054,
    input wire        mb1_FA1_TA1_IO_057_mb1_FB1_TA2_IO_055,
    input wire        mb1_FA1_TA1_IO_058_mb1_FB1_TA2_IO_072,
    input wire        mb1_FA1_TA1_IO_059_mb1_FB1_TA2_IO_073,
    input wire        mb1_FA1_TA1_IO_060_mb1_FB1_TA2_IO_070,
    input wire        mb1_FA1_TA1_IO_061_mb1_FB1_TA2_IO_071,
    input wire        mb1_FA1_TA1_IO_062_mb1_FB1_TA2_IO_048,
    input wire        mb1_FA1_TA1_IO_063_mb1_FB1_TA2_IO_049,
    input wire        mb1_FA1_TA1_IO_064_mb1_FB1_TA2_IO_066,
    input wire        mb1_FA1_TA1_IO_065_mb1_FB1_TA2_IO_067,
    input wire        mb1_FA1_TA1_IO_066_mb1_FB1_TA2_IO_064,
    input wire        mb1_FA1_TA1_IO_067_mb1_FB1_TA2_IO_065,
    input wire        mb1_FA1_TA1_IO_068_mb1_FB1_TA2_IO_082,
    input wire        mb1_FA1_TA1_IO_069_mb1_FB1_TA2_IO_083,
    input wire        mb1_FA1_TA1_IO_070_mb1_FB1_TA2_IO_060,
    input wire        mb1_FA1_TA1_IO_071_mb1_FB1_TA2_IO_061,
    input wire        mb1_FA1_TA1_IO_072_mb1_FB1_TA2_IO_058,
    input wire        mb1_FA1_TA1_IO_073_mb1_FB1_TA2_IO_059,
    input wire        mb1_FA1_TA1_IO_074_mb1_FB1_TA2_IO_076,
    input wire        mb1_FA1_TA1_IO_075_mb1_FB1_TA2_IO_077,
    input wire        mb1_FA1_TA1_IO_076_mb1_FB1_TA2_IO_074,
    input wire        mb1_FA1_TA1_IO_077_mb1_FB1_TA2_IO_075,
    input wire        mb1_FA1_TA1_IO_078_mb1_FB1_TA2_IO_092,
    input wire        mb1_FA1_TA1_IO_079_mb1_FB1_TA2_IO_093,
    input wire        mb1_FA1_TA1_IO_080_mb1_FB1_TA2_IO_090,
    input wire        mb1_FA1_TA1_IO_081_mb1_FB1_TA2_IO_091,
    input wire        mb1_FA1_TA1_IO_082_mb1_FB1_TA2_IO_068,
    input wire        mb1_FA1_TA1_IO_083_mb1_FB1_TA2_IO_069,
    input wire        mb1_FA1_TA1_IO_084_mb1_FB1_TA2_IO_086,
    input wire        mb1_FA1_TA1_IO_085_mb1_FB1_TA2_IO_087,
    input wire        mb1_FA1_TA1_IO_086_mb1_FB1_TA2_IO_084,
    input wire        mb1_FA1_TA1_IO_087_mb1_FB1_TA2_IO_085,
    input wire        mb1_FA1_TA1_IO_088_mb1_FB1_TA2_IO_102,
    input wire        mb1_FA1_TA1_IO_089_mb1_FB1_TA2_IO_103,
    input wire        mb1_FA1_TA1_IO_090_mb1_FB1_TA2_IO_080,
    input wire        mb1_FA1_TA1_IO_091_mb1_FB1_TA2_IO_081,
    input wire        mb1_FA1_TA1_IO_092_mb1_FB1_TA2_IO_078,
    input wire        mb1_FA1_TA1_IO_093_mb1_FB1_TA2_IO_079,
    input wire        mb1_FA1_TA1_IO_094_mb1_FB1_TA2_IO_096,
    input wire        mb1_FA1_TA1_IO_095_mb1_FB1_TA2_IO_097,
    input wire        mb1_FA1_TA1_IO_096_mb1_FB1_TA2_IO_094,
    input wire        mb1_FA1_TA1_IO_097_mb1_FB1_TA2_IO_095,
    input wire        mb1_FA1_TA1_IO_098_mb1_FB1_TA2_IO_112,
    input wire        mb1_FA1_TA1_IO_099_mb1_FB1_TA2_IO_113,
    input wire        mb1_FA1_TA1_IO_100_mb1_FB1_TA2_IO_110,
    input wire        mb1_FA1_TA1_IO_101_mb1_FB1_TA2_IO_111,
    input wire        mb1_FA1_TA1_IO_102_mb1_FB1_TA2_IO_088,
    input wire        mb1_FA1_TA1_IO_103_mb1_FB1_TA2_IO_089,
    input wire        mb1_FA1_TA1_IO_104_mb1_FB1_TA2_IO_106,
    input wire        mb1_FA1_TA1_IO_105_mb1_FB1_TA2_IO_107,
    input wire        mb1_FA1_TA1_IO_106_mb1_FB1_TA2_IO_104,
    input wire        mb1_FA1_TA1_IO_107_mb1_FB1_TA2_IO_105,
    input wire        mb1_FA1_TA1_IO_108_mb1_FB1_TA2_IO_122,
    input wire        mb1_FA1_TA1_IO_109_mb1_FB1_TA2_IO_123,
    input wire        mb1_FA1_TA1_IO_110_mb1_FB1_TA2_IO_100,
    input wire        mb1_FA1_TA1_IO_111_mb1_FB1_TA2_IO_101,
    input wire        mb1_FA1_TA1_IO_112_mb1_FB1_TA2_IO_098,
    input wire        mb1_FA1_TA1_IO_113_mb1_FB1_TA2_IO_099,
    input wire        mb1_FA1_TA1_IO_114_mb1_FB1_TA2_IO_116,
    input wire        mb1_FA1_TA1_IO_115_mb1_FB1_TA2_IO_117,
    input wire        mb1_FA1_TA1_IO_116_mb1_FB1_TA2_IO_114,
    input wire        mb1_FA1_TA1_IO_117_mb1_FB1_TA2_IO_115,
    input wire        mb1_FA1_TA1_IO_118_mb1_FB1_TA2_IO_132,
    input wire        mb1_FA1_TA1_IO_119_mb1_FB1_TA2_IO_133,
    input wire        mb1_FA1_TA1_IO_120_mb1_FB1_TA2_IO_130,
    input wire        mb1_FA1_TA1_IO_121_mb1_FB1_TA2_IO_131,
    input wire        mb1_FA1_TA1_IO_122_mb1_FB1_TA2_IO_108,
    input wire        mb1_FA1_TA1_IO_123_mb1_FB1_TA2_IO_109,
    input wire        mb1_FA1_TA1_IO_124_mb1_FB1_TA2_IO_126,
    input wire        mb1_FA1_TA1_IO_125_mb1_FB1_TA2_IO_127,
    input wire        mb1_FA1_TA1_IO_126_mb1_FB1_TA2_IO_124,
    input wire        mb1_FA1_TA1_IO_127_mb1_FB1_TA2_IO_125,
    input wire        mb1_FA1_TA1_IO_130_mb1_FB1_TA2_IO_120,
    input wire        mb1_FA1_TA1_IO_131_mb1_FB1_TA2_IO_121,
    input wire        mb1_FA1_TA1_IO_132_mb1_FB1_TA2_IO_118,
    input wire        mb1_FA1_TA1_IO_133_mb1_FB1_TA2_IO_119,
    input wire        mb1_FA1_TA1_IO_134_mb1_FB1_TA2_IO_136,
    input wire        mb1_FA1_TA1_IO_136_mb1_FB1_TA2_IO_134,
    output wire        mb1_FB1_TB0_CLKIO_N_0_mb1_FB2_BB2_CLKIO_N_7,
    output wire        mb1_FB1_TB0_CLKIO_N_1_mb1_FB2_BB2_CLKIO_N_6,
    output wire        mb1_FB1_TB0_CLKIO_N_2_mb1_FB2_BB2_CLKIO_N_4,
    output wire        mb1_FB1_TB0_CLKIO_N_3_mb1_FB2_BB2_CLKIO_N_3,
    output wire        mb1_FB1_TB0_CLKIO_N_4_mb1_FB2_BB2_CLKIO_N_2,
    output wire        mb1_FB1_TB0_CLKIO_N_5_mb1_FB2_BB2_IO_010,
    output wire        mb1_FB1_TB0_CLKIO_N_6_mb1_FB2_BB2_CLKIO_N_1,
    output wire        mb1_FB1_TB0_CLKIO_N_7_mb1_FB2_BB2_CLKIO_N_0,
    output wire        mb1_FB1_TB0_CLKIO_P_0_mb1_FB2_BB2_CLKIO_P_7,
    output wire        mb1_FB1_TB0_CLKIO_P_1_mb1_FB2_BB2_CLKIO_P_6,
    output wire        mb1_FB1_TB0_CLKIO_P_2_mb1_FB2_BB2_CLKIO_P_4,
    output wire        mb1_FB1_TB0_CLKIO_P_3_mb1_FB2_BB2_CLKIO_P_3,
    output wire        mb1_FB1_TB0_CLKIO_P_4_mb1_FB2_BB2_CLKIO_P_2,
    output wire        mb1_FB1_TB0_CLKIO_P_5_mb1_FB2_BB2_IO_011,
    output wire        mb1_FB1_TB0_CLKIO_P_6_mb1_FB2_BB2_CLKIO_P_1,
    output wire        mb1_FB1_TB0_CLKIO_P_7_mb1_FB2_BB2_CLKIO_P_0,
    output wire        mb1_FB1_TB0_IO_004_mb1_FB2_BB2_IO_006,
    output wire        mb1_FB1_TB0_IO_005_mb1_FB2_BB2_IO_007,
    output wire        mb1_FB1_TB0_IO_006_mb1_FB2_BB2_IO_004,
    output wire        mb1_FB1_TB0_IO_007_mb1_FB2_BB2_IO_005,
    output wire        mb1_FB1_TB0_IO_008_mb1_FB2_BB2_IO_022,
    output wire        mb1_FB1_TB0_IO_009_mb1_FB2_BB2_IO_023,
    output wire        mb1_FB1_TB0_IO_010_mb1_FB2_BB2_CLKIO_N_5,
    output wire        mb1_FB1_TB0_IO_011_mb1_FB2_BB2_CLKIO_P_5,
    output wire        mb1_FB1_TB0_IO_012_mb1_FB2_BB2_IO_012,
    output wire        mb1_FB1_TB0_IO_013_mb1_FB2_BB2_IO_013,
    output wire        mb1_FB1_TB0_IO_014_mb1_FB2_BB2_IO_016,
    output wire        mb1_FB1_TB0_IO_015_mb1_FB2_BB2_IO_017,
    output wire        mb1_FB1_TB0_IO_016_mb1_FB2_BB2_IO_014,
    output wire        mb1_FB1_TB0_IO_017_mb1_FB2_BB2_IO_015,
    output wire        mb1_FB1_TB0_IO_018_mb1_FB2_BB2_IO_032,
    output wire        mb1_FB1_TB0_IO_019_mb1_FB2_BB2_IO_033,
    output wire        mb1_FB1_TB0_IO_020_mb1_FB2_BB2_IO_030,
    output wire        mb1_FB1_TB0_IO_021_mb1_FB2_BB2_IO_031,
    output wire        mb1_FB1_TB0_IO_022_mb1_FB2_BB2_IO_008,
    output wire        mb1_FB1_TB0_IO_023_mb1_FB2_BB2_IO_009,
    output wire        mb1_FB1_TB0_IO_024_mb1_FB2_BB2_IO_026,
    output wire        mb1_FB1_TB0_IO_025_mb1_FB2_BB2_IO_027,
    output wire        mb1_FB1_TB0_IO_026_mb1_FB2_BB2_IO_024,
    output wire        mb1_FB1_TB0_IO_027_mb1_FB2_BB2_IO_025,
    output wire        mb1_FB1_TB0_IO_028_mb1_FB2_BB2_IO_042,
    output wire        mb1_FB1_TB0_IO_029_mb1_FB2_BB2_IO_043,
    output wire        mb1_FB1_TB0_IO_030_mb1_FB2_BB2_IO_020,
    output wire        mb1_FB1_TB0_IO_031_mb1_FB2_BB2_IO_021,
    output wire        mb1_FB1_TB0_IO_032_mb1_FB2_BB2_IO_018,
    output wire        mb1_FB1_TB0_IO_033_mb1_FB2_BB2_IO_019,
    output wire        mb1_FB1_TB0_IO_034_mb1_FB2_BB2_IO_036,
    output wire        mb1_FB1_TB0_IO_035_mb1_FB2_BB2_IO_037,
    output wire        mb1_FB1_TB0_IO_036_mb1_FB2_BB2_IO_034,
    output wire        mb1_FB1_TB0_IO_037_mb1_FB2_BB2_IO_035,
    output wire        mb1_FB1_TB0_IO_038_mb1_FB2_BB2_IO_052,
    output wire        mb1_FB1_TB0_IO_039_mb1_FB2_BB2_IO_053,
    output wire        mb1_FB1_TB0_IO_040_mb1_FB2_BB2_IO_050,
    output wire        mb1_FB1_TB0_IO_041_mb1_FB2_BB2_IO_051,
    output wire        mb1_FB1_TB0_IO_042_mb1_FB2_BB2_IO_028,
    output wire        mb1_FB1_TB0_IO_043_mb1_FB2_BB2_IO_029,
    output wire        mb1_FB1_TB0_IO_044_mb1_FB2_BB2_IO_046,
    output wire        mb1_FB1_TB0_IO_045_mb1_FB2_BB2_IO_047,
    output wire        mb1_FB1_TB0_IO_046_mb1_FB2_BB2_IO_044,
    output wire        mb1_FB1_TB0_IO_047_mb1_FB2_BB2_IO_045,
    output wire        mb1_FB1_TB0_IO_048_mb1_FB2_BB2_IO_062,
    output wire        mb1_FB1_TB0_IO_049_mb1_FB2_BB2_IO_063,
    output wire        mb1_FB1_TB0_IO_050_mb1_FB2_BB2_IO_040,
    output wire        mb1_FB1_TB0_IO_051_mb1_FB2_BB2_IO_041,
    output wire        mb1_FB1_TB0_IO_052_mb1_FB2_BB2_IO_038,
    output wire        mb1_FB1_TB0_IO_053_mb1_FB2_BB2_IO_039,
    output wire        mb1_FB1_TB0_IO_054_mb1_FB2_BB2_IO_056,
    output wire        mb1_FB1_TB0_IO_055_mb1_FB2_BB2_IO_057,
    output wire        mb1_FB1_TB0_IO_056_mb1_FB2_BB2_IO_054,
    output wire        mb1_FB1_TB0_IO_057_mb1_FB2_BB2_IO_055,
    output wire        mb1_FB1_TB0_IO_058_mb1_FB2_BB2_IO_072,
    output wire        mb1_FB1_TB0_IO_059_mb1_FB2_BB2_IO_073,
    output wire        mb1_FB1_TB0_IO_060_mb1_FB2_BB2_IO_070,
    output wire        mb1_FB1_TB0_IO_061_mb1_FB2_BB2_IO_071,
    output wire        mb1_FB1_TB0_IO_062_mb1_FB2_BB2_IO_048,
    output wire        mb1_FB1_TB0_IO_063_mb1_FB2_BB2_IO_049,
    output wire        mb1_FB1_TB0_IO_064_mb1_FB2_BB2_IO_066,
    output wire        mb1_FB1_TB0_IO_065_mb1_FB2_BB2_IO_067,
    output wire        mb1_FB1_TB0_IO_066_mb1_FB2_BB2_IO_064,
    output wire        mb1_FB1_TB0_IO_067_mb1_FB2_BB2_IO_065,
    output wire        mb1_FB1_TB0_IO_068_mb1_FB2_BB2_IO_082,
    output wire        mb1_FB1_TB0_IO_069_mb1_FB2_BB2_IO_083,
    output wire        mb1_FB1_TB0_IO_070_mb1_FB2_BB2_IO_060,
    output wire        mb1_FB1_TB0_IO_071_mb1_FB2_BB2_IO_061,
    output wire        mb1_FB1_TB0_IO_072_mb1_FB2_BB2_IO_058,
    output wire        mb1_FB1_TB0_IO_073_mb1_FB2_BB2_IO_059,
    output wire        mb1_FB1_TB0_IO_074_mb1_FB2_BB2_IO_076,
    output wire        mb1_FB1_TB0_IO_075_mb1_FB2_BB2_IO_077,
    output wire        mb1_FB1_TB0_IO_076_mb1_FB2_BB2_IO_074,
    output wire        mb1_FB1_TB0_IO_077_mb1_FB2_BB2_IO_075,
    output wire        mb1_FB1_TB0_IO_078_mb1_FB2_BB2_IO_092,
    output wire        mb1_FB1_TB0_IO_079_mb1_FB2_BB2_IO_093,
    output wire        mb1_FB1_TB0_IO_080_mb1_FB2_BB2_IO_090,
    output wire        mb1_FB1_TB0_IO_081_mb1_FB2_BB2_IO_091,
    output wire        mb1_FB1_TB0_IO_082_mb1_FB2_BB2_IO_068,
    output wire        mb1_FB1_TB0_IO_083_mb1_FB2_BB2_IO_069,
    output wire        mb1_FB1_TB0_IO_084_mb1_FB2_BB2_IO_086,
    output wire        mb1_FB1_TB0_IO_085_mb1_FB2_BB2_IO_087,
    output wire        mb1_FB1_TB0_IO_086_mb1_FB2_BB2_IO_084,
    output wire        mb1_FB1_TB0_IO_087_mb1_FB2_BB2_IO_085,
    output wire        mb1_FB1_TB0_IO_088_mb1_FB2_BB2_IO_102,
    output wire        mb1_FB1_TB0_IO_089_mb1_FB2_BB2_IO_103,
    output wire        mb1_FB1_TB0_IO_090_mb1_FB2_BB2_IO_080,
    output wire        mb1_FB1_TB0_IO_091_mb1_FB2_BB2_IO_081,
    output wire        mb1_FB1_TB0_IO_092_mb1_FB2_BB2_IO_078,
    output wire        mb1_FB1_TB0_IO_093_mb1_FB2_BB2_IO_079,
    output wire        mb1_FB1_TB0_IO_094_mb1_FB2_BB2_IO_096,
    output wire        mb1_FB1_TB0_IO_095_mb1_FB2_BB2_IO_097,
    output wire        mb1_FB1_TB0_IO_096_mb1_FB2_BB2_IO_094,
    output wire        mb1_FB1_TB0_IO_097_mb1_FB2_BB2_IO_095,
    output wire        mb1_FB1_TB0_IO_098_mb1_FB2_BB2_IO_112,
    output wire        mb1_FB1_TB0_IO_099_mb1_FB2_BB2_IO_113,
    output wire        mb1_FB1_TB0_IO_100_mb1_FB2_BB2_IO_110,
    output wire        mb1_FB1_TB0_IO_101_mb1_FB2_BB2_IO_111,
    output wire        mb1_FB1_TB0_IO_102_mb1_FB2_BB2_IO_088,
    output wire        mb1_FB1_TB0_IO_103_mb1_FB2_BB2_IO_089,
    output wire        mb1_FB1_TB0_IO_104_mb1_FB2_BB2_IO_106,
    output wire        mb1_FB1_TB0_IO_105_mb1_FB2_BB2_IO_107,
    output wire        mb1_FB1_TB0_IO_106_mb1_FB2_BB2_IO_104,
    output wire        mb1_FB1_TB0_IO_107_mb1_FB2_BB2_IO_105,
    output wire        mb1_FB1_TB0_IO_108_mb1_FB2_BB2_IO_122,
    output wire        mb1_FB1_TB0_IO_109_mb1_FB2_BB2_IO_123,
    output wire        mb1_FB1_TB0_IO_110_mb1_FB2_BB2_IO_100,
    output wire        mb1_FB1_TB0_IO_111_mb1_FB2_BB2_IO_101,
    output wire        mb1_FB1_TB0_IO_112_mb1_FB2_BB2_IO_098,
    output wire        mb1_FB1_TB0_IO_113_mb1_FB2_BB2_IO_099,
    output wire        mb1_FB1_TB0_IO_114_mb1_FB2_BB2_IO_116,
    output wire        mb1_FB1_TB0_IO_115_mb1_FB2_BB2_IO_117,
    output wire        mb1_FB1_TB0_IO_116_mb1_FB2_BB2_IO_114,
    output wire        mb1_FB1_TB0_IO_117_mb1_FB2_BB2_IO_115,
    output wire        mb1_FB1_TB0_IO_118_mb1_FB2_BB2_IO_132,
    output wire        mb1_FB1_TB0_IO_119_mb1_FB2_BB2_IO_133,
    output wire        mb1_FB1_TB0_IO_120_mb1_FB2_BB2_IO_130,
    output wire        mb1_FB1_TB0_IO_121_mb1_FB2_BB2_IO_131,
    output wire        mb1_FB1_TB0_IO_122_mb1_FB2_BB2_IO_108,
    output wire        mb1_FB1_TB0_IO_123_mb1_FB2_BB2_IO_109,
    output wire        mb1_FB1_TB0_IO_124_mb1_FB2_BB2_IO_126,
    output wire        mb1_FB1_TB0_IO_125_mb1_FB2_BB2_IO_127,
    output wire        mb1_FB1_TB0_IO_126_mb1_FB2_BB2_IO_124,
    output wire        mb1_FB1_TB0_IO_127_mb1_FB2_BB2_IO_125,
    output wire        mb1_FB1_TB0_IO_130_mb1_FB2_BB2_IO_120,
    output wire        mb1_FB1_TB0_IO_131_mb1_FB2_BB2_IO_121,
    output wire        mb1_FB1_TB0_IO_132_mb1_FB2_BB2_IO_118,
    output wire        mb1_FB1_TB0_IO_133_mb1_FB2_BB2_IO_119,
    output wire        mb1_FB1_TB0_IO_134_mb1_FB2_BB2_IO_136,
    output wire        mb1_FB1_TB0_IO_136_mb1_FB2_BB2_IO_134,
    output wire        mb1_FB1_TB1_CLKIO_N_0_mb1_FA2_BA1_CLKIO_N_7,
    output wire        mb1_FB1_TB1_CLKIO_N_1_mb1_FA2_BA1_CLKIO_N_6,
    output wire        mb1_FB1_TB1_CLKIO_N_2_mb1_FA2_BA1_CLKIO_N_4,
    output wire        mb1_FB1_TB1_CLKIO_N_3_mb1_FA2_BA1_CLKIO_N_3,
    output wire        mb1_FB1_TB1_CLKIO_N_4_mb1_FA2_BA1_CLKIO_N_2,
    output wire        mb1_FB1_TB1_CLKIO_N_5_mb1_FA2_BA1_IO_010,
    output wire        mb1_FB1_TB1_CLKIO_N_6_mb1_FA2_BA1_CLKIO_N_1,
    output wire        mb1_FB1_TB1_CLKIO_N_7_mb1_FA2_BA1_CLKIO_N_0,
    output wire        mb1_FB1_TB1_CLKIO_P_0_mb1_FA2_BA1_CLKIO_P_7,
    output wire        mb1_FB1_TB1_CLKIO_P_1_mb1_FA2_BA1_CLKIO_P_6,
    output wire        mb1_FB1_TB1_CLKIO_P_2_mb1_FA2_BA1_CLKIO_P_4,
    output wire        mb1_FB1_TB1_CLKIO_P_3_mb1_FA2_BA1_CLKIO_P_3,
    output wire        mb1_FB1_TB1_CLKIO_P_4_mb1_FA2_BA1_CLKIO_P_2,
    output wire        mb1_FB1_TB1_CLKIO_P_5_mb1_FA2_BA1_IO_011,
    output wire        mb1_FB1_TB1_CLKIO_P_6_mb1_FA2_BA1_CLKIO_P_1,
    output wire        mb1_FB1_TB1_CLKIO_P_7_mb1_FA2_BA1_CLKIO_P_0,
    output wire        mb1_FB1_TB1_IO_004_mb1_FA2_BA1_IO_006,
    output wire        mb1_FB1_TB1_IO_005_mb1_FA2_BA1_IO_007,
    output wire        mb1_FB1_TB1_IO_006_mb1_FA2_BA1_IO_004,
    output wire        mb1_FB1_TB1_IO_007_mb1_FA2_BA1_IO_005,
    output wire        mb1_FB1_TB1_IO_008_mb1_FA2_BA1_IO_022,
    output wire        mb1_FB1_TB1_IO_009_mb1_FA2_BA1_IO_023,
    output wire        mb1_FB1_TB1_IO_010_mb1_FA2_BA1_CLKIO_N_5,
    output wire        mb1_FB1_TB1_IO_011_mb1_FA2_BA1_CLKIO_P_5,
    output wire        mb1_FB1_TB1_IO_012_mb1_FA2_BA1_IO_012,
    output wire        mb1_FB1_TB1_IO_013_mb1_FA2_BA1_IO_013,
    output wire        mb1_FB1_TB1_IO_014_mb1_FA2_BA1_IO_016,
    output wire        mb1_FB1_TB1_IO_015_mb1_FA2_BA1_IO_017,
    output wire        mb1_FB1_TB1_IO_016_mb1_FA2_BA1_IO_014,
    output wire        mb1_FB1_TB1_IO_017_mb1_FA2_BA1_IO_015,
    output wire        mb1_FB1_TB1_IO_018_mb1_FA2_BA1_IO_032,
    output wire        mb1_FB1_TB1_IO_019_mb1_FA2_BA1_IO_033,
    output wire        mb1_FB1_TB1_IO_020_mb1_FA2_BA1_IO_030,
    output wire        mb1_FB1_TB1_IO_021_mb1_FA2_BA1_IO_031,
    output wire        mb1_FB1_TB1_IO_022_mb1_FA2_BA1_IO_008,
    output wire        mb1_FB1_TB1_IO_023_mb1_FA2_BA1_IO_009,
    output wire        mb1_FB1_TB1_IO_024_mb1_FA2_BA1_IO_026,
    output wire        mb1_FB1_TB1_IO_025_mb1_FA2_BA1_IO_027,
    output wire        mb1_FB1_TB1_IO_026_mb1_FA2_BA1_IO_024,
    output wire        mb1_FB1_TB1_IO_027_mb1_FA2_BA1_IO_025,
    output wire        mb1_FB1_TB1_IO_028_mb1_FA2_BA1_IO_042,
    output wire        mb1_FB1_TB1_IO_029_mb1_FA2_BA1_IO_043,
    output wire        mb1_FB1_TB1_IO_030_mb1_FA2_BA1_IO_020,
    output wire        mb1_FB1_TB1_IO_031_mb1_FA2_BA1_IO_021,
    output wire        mb1_FB1_TB1_IO_032_mb1_FA2_BA1_IO_018,
    output wire        mb1_FB1_TB1_IO_033_mb1_FA2_BA1_IO_019,
    output wire        mb1_FB1_TB1_IO_034_mb1_FA2_BA1_IO_036,
    output wire        mb1_FB1_TB1_IO_035_mb1_FA2_BA1_IO_037,
    output wire        mb1_FB1_TB1_IO_036_mb1_FA2_BA1_IO_034,
    output wire        mb1_FB1_TB1_IO_037_mb1_FA2_BA1_IO_035,
    output wire        mb1_FB1_TB1_IO_038_mb1_FA2_BA1_IO_052,
    output wire        mb1_FB1_TB1_IO_039_mb1_FA2_BA1_IO_053,
    output wire        mb1_FB1_TB1_IO_040_mb1_FA2_BA1_IO_050,
    output wire        mb1_FB1_TB1_IO_041_mb1_FA2_BA1_IO_051,
    output wire        mb1_FB1_TB1_IO_042_mb1_FA2_BA1_IO_028,
    output wire        mb1_FB1_TB1_IO_043_mb1_FA2_BA1_IO_029,
    output wire        mb1_FB1_TB1_IO_044_mb1_FA2_BA1_IO_046,
    output wire        mb1_FB1_TB1_IO_045_mb1_FA2_BA1_IO_047,
    output wire        mb1_FB1_TB1_IO_046_mb1_FA2_BA1_IO_044,
    output wire        mb1_FB1_TB1_IO_047_mb1_FA2_BA1_IO_045,
    output wire        mb1_FB1_TB1_IO_048_mb1_FA2_BA1_IO_062,
    output wire        mb1_FB1_TB1_IO_049_mb1_FA2_BA1_IO_063,
    output wire        mb1_FB1_TB1_IO_050_mb1_FA2_BA1_IO_040,
    output wire        mb1_FB1_TB1_IO_051_mb1_FA2_BA1_IO_041,
    output wire        mb1_FB1_TB1_IO_052_mb1_FA2_BA1_IO_038,
    output wire        mb1_FB1_TB1_IO_053_mb1_FA2_BA1_IO_039,
    output wire        mb1_FB1_TB1_IO_054_mb1_FA2_BA1_IO_056,
    output wire        mb1_FB1_TB1_IO_055_mb1_FA2_BA1_IO_057,
    output wire        mb1_FB1_TB1_IO_056_mb1_FA2_BA1_IO_054,
    output wire        mb1_FB1_TB1_IO_057_mb1_FA2_BA1_IO_055,
    output wire        mb1_FB1_TB1_IO_058_mb1_FA2_BA1_IO_072,
    output wire        mb1_FB1_TB1_IO_059_mb1_FA2_BA1_IO_073,
    output wire        mb1_FB1_TB1_IO_060_mb1_FA2_BA1_IO_070,
    output wire        mb1_FB1_TB1_IO_061_mb1_FA2_BA1_IO_071,
    output wire        mb1_FB1_TB1_IO_062_mb1_FA2_BA1_IO_048,
    output wire        mb1_FB1_TB1_IO_063_mb1_FA2_BA1_IO_049,
    output wire        mb1_FB1_TB1_IO_064_mb1_FA2_BA1_IO_066,
    output wire        mb1_FB1_TB1_IO_065_mb1_FA2_BA1_IO_067,
    output wire        mb1_FB1_TB1_IO_066_mb1_FA2_BA1_IO_064,
    output wire        mb1_FB1_TB1_IO_067_mb1_FA2_BA1_IO_065,
    output wire        mb1_FB1_TB1_IO_068_mb1_FA2_BA1_IO_082,
    output wire        mb1_FB1_TB1_IO_069_mb1_FA2_BA1_IO_083,
    output wire        mb1_FB1_TB1_IO_070_mb1_FA2_BA1_IO_060,
    output wire        mb1_FB1_TB1_IO_071_mb1_FA2_BA1_IO_061,
    output wire        mb1_FB1_TB1_IO_072_mb1_FA2_BA1_IO_058,
    output wire        mb1_FB1_TB1_IO_073_mb1_FA2_BA1_IO_059,
    output wire        mb1_FB1_TB1_IO_074_mb1_FA2_BA1_IO_076,
    output wire        mb1_FB1_TB1_IO_075_mb1_FA2_BA1_IO_077,
    output wire        mb1_FB1_TB1_IO_076_mb1_FA2_BA1_IO_074,
    output wire        mb1_FB1_TB1_IO_077_mb1_FA2_BA1_IO_075,
    output wire        mb1_FB1_TB1_IO_078_mb1_FA2_BA1_IO_092,
    output wire        mb1_FB1_TB1_IO_079_mb1_FA2_BA1_IO_093,
    output wire        mb1_FB1_TB1_IO_080_mb1_FA2_BA1_IO_090,
    output wire        mb1_FB1_TB1_IO_081_mb1_FA2_BA1_IO_091,
    output wire        mb1_FB1_TB1_IO_082_mb1_FA2_BA1_IO_068,
    output wire        mb1_FB1_TB1_IO_083_mb1_FA2_BA1_IO_069,
    output wire        mb1_FB1_TB1_IO_084_mb1_FA2_BA1_IO_086,
    output wire        mb1_FB1_TB1_IO_085_mb1_FA2_BA1_IO_087,
    output wire        mb1_FB1_TB1_IO_086_mb1_FA2_BA1_IO_084,
    output wire        mb1_FB1_TB1_IO_087_mb1_FA2_BA1_IO_085,
    output wire        mb1_FB1_TB1_IO_088_mb1_FA2_BA1_IO_102,
    output wire        mb1_FB1_TB1_IO_089_mb1_FA2_BA1_IO_103,
    output wire        mb1_FB1_TB1_IO_090_mb1_FA2_BA1_IO_080,
    output wire        mb1_FB1_TB1_IO_091_mb1_FA2_BA1_IO_081,
    output wire        mb1_FB1_TB1_IO_092_mb1_FA2_BA1_IO_078,
    output wire        mb1_FB1_TB1_IO_093_mb1_FA2_BA1_IO_079,
    output wire        mb1_FB1_TB1_IO_094_mb1_FA2_BA1_IO_096,
    output wire        mb1_FB1_TB1_IO_095_mb1_FA2_BA1_IO_097,
    output wire        mb1_FB1_TB1_IO_096_mb1_FA2_BA1_IO_094,
    output wire        mb1_FB1_TB1_IO_097_mb1_FA2_BA1_IO_095,
    output wire        mb1_FB1_TB1_IO_098_mb1_FA2_BA1_IO_112,
    output wire        mb1_FB1_TB1_IO_099_mb1_FA2_BA1_IO_113,
    output wire        mb1_FB1_TB1_IO_100_mb1_FA2_BA1_IO_110,
    output wire        mb1_FB1_TB1_IO_101_mb1_FA2_BA1_IO_111,
    output wire        mb1_FB1_TB1_IO_102_mb1_FA2_BA1_IO_088,
    output wire        mb1_FB1_TB1_IO_103_mb1_FA2_BA1_IO_089,
    output wire        mb1_FB1_TB1_IO_104_mb1_FA2_BA1_IO_106,
    output wire        mb1_FB1_TB1_IO_105_mb1_FA2_BA1_IO_107,
    output wire        mb1_FB1_TB1_IO_106_mb1_FA2_BA1_IO_104,
    output wire        mb1_FB1_TB1_IO_107_mb1_FA2_BA1_IO_105,
    output wire        mb1_FB1_TB1_IO_108_mb1_FA2_BA1_IO_122,
    output wire        mb1_FB1_TB1_IO_109_mb1_FA2_BA1_IO_123,
    output wire        mb1_FB1_TB1_IO_110_mb1_FA2_BA1_IO_100,
    output wire        mb1_FB1_TB1_IO_111_mb1_FA2_BA1_IO_101,
    output wire        mb1_FB1_TB1_IO_112_mb1_FA2_BA1_IO_098,
    output wire        mb1_FB1_TB1_IO_113_mb1_FA2_BA1_IO_099,
    output wire        mb1_FB1_TB1_IO_114_mb1_FA2_BA1_IO_116,
    output wire        mb1_FB1_TB1_IO_115_mb1_FA2_BA1_IO_117,
    output wire        mb1_FB1_TB1_IO_116_mb1_FA2_BA1_IO_114,
    output wire        mb1_FB1_TB1_IO_117_mb1_FA2_BA1_IO_115,
    output wire        mb1_FB1_TB1_IO_118_mb1_FA2_BA1_IO_132,
    output wire        mb1_FB1_TB1_IO_119_mb1_FA2_BA1_IO_133,
    output wire        mb1_FB1_TB1_IO_120_mb1_FA2_BA1_IO_130,
    output wire        mb1_FB1_TB1_IO_121_mb1_FA2_BA1_IO_131,
    output wire        mb1_FB1_TB1_IO_122_mb1_FA2_BA1_IO_108,
    output wire        mb1_FB1_TB1_IO_123_mb1_FA2_BA1_IO_109,
    output wire        mb1_FB1_TB1_IO_124_mb1_FA2_BA1_IO_126,
    output wire        mb1_FB1_TB1_IO_125_mb1_FA2_BA1_IO_127,
    output wire        mb1_FB1_TB1_IO_126_mb1_FA2_BA1_IO_124,
    output wire        mb1_FB1_TB1_IO_127_mb1_FA2_BA1_IO_125,
    output wire        mb1_FB1_TB1_IO_130_mb1_FA2_BA1_IO_120,
    output wire        mb1_FB1_TB1_IO_131_mb1_FA2_BA1_IO_121,
    output wire        mb1_FB1_TB1_IO_132_mb1_FA2_BA1_IO_118,
    output wire        mb1_FB1_TB1_IO_133_mb1_FA2_BA1_IO_119,
    output wire        mb1_FB1_TB1_IO_134_mb1_FA2_BA1_IO_136,
    output wire        mb1_FB1_TB1_IO_136_mb1_FA2_BA1_IO_134,
    input wire        mb1_FA1_TB0_CLKIO_N_0_mb1_FB1_TB2_CLKIO_N_7,
    input wire        mb1_FA1_TB0_CLKIO_N_1_mb1_FB1_TB2_CLKIO_N_6,
    input wire        mb1_FA1_TB0_CLKIO_N_2_mb1_FB1_TB2_CLKIO_N_4,
    input wire        mb1_FA1_TB0_CLKIO_N_3_mb1_FB1_TB2_CLKIO_N_3,
    input wire        mb1_FA1_TB0_CLKIO_N_4_mb1_FB1_TB2_CLKIO_N_2,
    input wire        mb1_FA1_TB0_CLKIO_N_5_mb1_FB1_TB2_IO_010,
    input wire        mb1_FA1_TB0_CLKIO_N_6_mb1_FB1_TB2_CLKIO_N_1,
    input wire        mb1_FA1_TB0_CLKIO_N_7_mb1_FB1_TB2_CLKIO_N_0,
    input wire        mb1_FA1_TB0_CLKIO_P_0_mb1_FB1_TB2_CLKIO_P_7,
    input wire        mb1_FA1_TB0_CLKIO_P_1_mb1_FB1_TB2_CLKIO_P_6,
    input wire        mb1_FA1_TB0_CLKIO_P_2_mb1_FB1_TB2_CLKIO_P_4,
    input wire        mb1_FA1_TB0_CLKIO_P_3_mb1_FB1_TB2_CLKIO_P_3,
    input wire        mb1_FA1_TB0_CLKIO_P_4_mb1_FB1_TB2_CLKIO_P_2,
    input wire        mb1_FA1_TB0_CLKIO_P_5_mb1_FB1_TB2_IO_011,
    input wire        mb1_FA1_TB0_CLKIO_P_6_mb1_FB1_TB2_CLKIO_P_1,
    input wire        mb1_FA1_TB0_CLKIO_P_7_mb1_FB1_TB2_CLKIO_P_0,
    input wire        mb1_FA1_TB0_IO_004_mb1_FB1_TB2_IO_006,
    input wire        mb1_FA1_TB0_IO_005_mb1_FB1_TB2_IO_007,
    input wire        mb1_FA1_TB0_IO_006_mb1_FB1_TB2_IO_004,
    input wire        mb1_FA1_TB0_IO_007_mb1_FB1_TB2_IO_005,
    input wire        mb1_FA1_TB0_IO_008_mb1_FB1_TB2_IO_022,
    input wire        mb1_FA1_TB0_IO_009_mb1_FB1_TB2_IO_023,
    input wire        mb1_FA1_TB0_IO_010_mb1_FB1_TB2_CLKIO_N_5,
    input wire        mb1_FA1_TB0_IO_011_mb1_FB1_TB2_CLKIO_P_5,
    input wire        mb1_FA1_TB0_IO_012_mb1_FB1_TB2_IO_012,
    input wire        mb1_FA1_TB0_IO_013_mb1_FB1_TB2_IO_013,
    input wire        mb1_FA1_TB0_IO_014_mb1_FB1_TB2_IO_016,
    input wire        mb1_FA1_TB0_IO_015_mb1_FB1_TB2_IO_017,
    input wire        mb1_FA1_TB0_IO_016_mb1_FB1_TB2_IO_014,
    input wire        mb1_FA1_TB0_IO_017_mb1_FB1_TB2_IO_015,
    input wire        mb1_FA1_TB0_IO_018_mb1_FB1_TB2_IO_032,
    input wire        mb1_FA1_TB0_IO_019_mb1_FB1_TB2_IO_033,
    input wire        mb1_FA1_TB0_IO_020_mb1_FB1_TB2_IO_030,
    input wire        mb1_FA1_TB0_IO_021_mb1_FB1_TB2_IO_031,
    input wire        mb1_FA1_TB0_IO_022_mb1_FB1_TB2_IO_008,
    input wire        mb1_FA1_TB0_IO_023_mb1_FB1_TB2_IO_009,
    input wire        mb1_FA1_TB0_IO_024_mb1_FB1_TB2_IO_026,
    input wire        mb1_FA1_TB0_IO_025_mb1_FB1_TB2_IO_027,
    input wire        mb1_FA1_TB0_IO_026_mb1_FB1_TB2_IO_024,
    input wire        mb1_FA1_TB0_IO_027_mb1_FB1_TB2_IO_025,
    input wire        mb1_FA1_TB0_IO_028_mb1_FB1_TB2_IO_042,
    input wire        mb1_FA1_TB0_IO_029_mb1_FB1_TB2_IO_043,
    input wire        mb1_FA1_TB0_IO_030_mb1_FB1_TB2_IO_020,
    input wire        mb1_FA1_TB0_IO_031_mb1_FB1_TB2_IO_021,
    input wire        mb1_FA1_TB0_IO_032_mb1_FB1_TB2_IO_018,
    input wire        mb1_FA1_TB0_IO_033_mb1_FB1_TB2_IO_019,
    input wire        mb1_FA1_TB0_IO_034_mb1_FB1_TB2_IO_036,
    input wire        mb1_FA1_TB0_IO_035_mb1_FB1_TB2_IO_037,
    input wire        mb1_FA1_TB0_IO_036_mb1_FB1_TB2_IO_034,
    input wire        mb1_FA1_TB0_IO_037_mb1_FB1_TB2_IO_035,
    input wire        mb1_FA1_TB0_IO_038_mb1_FB1_TB2_IO_052,
    input wire        mb1_FA1_TB0_IO_039_mb1_FB1_TB2_IO_053,
    input wire        mb1_FA1_TB0_IO_040_mb1_FB1_TB2_IO_050,
    input wire        mb1_FA1_TB0_IO_041_mb1_FB1_TB2_IO_051,
    input wire        mb1_FA1_TB0_IO_042_mb1_FB1_TB2_IO_028,
    input wire        mb1_FA1_TB0_IO_043_mb1_FB1_TB2_IO_029,
    input wire        mb1_FA1_TB0_IO_044_mb1_FB1_TB2_IO_046,
    input wire        mb1_FA1_TB0_IO_045_mb1_FB1_TB2_IO_047,
    input wire        mb1_FA1_TB0_IO_046_mb1_FB1_TB2_IO_044,
    input wire        mb1_FA1_TB0_IO_047_mb1_FB1_TB2_IO_045,
    input wire        mb1_FA1_TB0_IO_048_mb1_FB1_TB2_IO_062,
    input wire        mb1_FA1_TB0_IO_049_mb1_FB1_TB2_IO_063,
    input wire        mb1_FA1_TB0_IO_050_mb1_FB1_TB2_IO_040,
    input wire        mb1_FA1_TB0_IO_051_mb1_FB1_TB2_IO_041,
    input wire        mb1_FA1_TB0_IO_052_mb1_FB1_TB2_IO_038,
    input wire        mb1_FA1_TB0_IO_053_mb1_FB1_TB2_IO_039,
    input wire        mb1_FA1_TB0_IO_054_mb1_FB1_TB2_IO_056,
    input wire        mb1_FA1_TB0_IO_055_mb1_FB1_TB2_IO_057,
    input wire        mb1_FA1_TB0_IO_056_mb1_FB1_TB2_IO_054,
    input wire        mb1_FA1_TB0_IO_057_mb1_FB1_TB2_IO_055,
    input wire        mb1_FA1_TB0_IO_058_mb1_FB1_TB2_IO_072,
    input wire        mb1_FA1_TB0_IO_059_mb1_FB1_TB2_IO_073,
    input wire        mb1_FA1_TB0_IO_060_mb1_FB1_TB2_IO_070,
    input wire        mb1_FA1_TB0_IO_061_mb1_FB1_TB2_IO_071,
    input wire        mb1_FA1_TB0_IO_062_mb1_FB1_TB2_IO_048,
    input wire        mb1_FA1_TB0_IO_063_mb1_FB1_TB2_IO_049,
    input wire        mb1_FA1_TB0_IO_064_mb1_FB1_TB2_IO_066,
    input wire        mb1_FA1_TB0_IO_065_mb1_FB1_TB2_IO_067,
    input wire        mb1_FA1_TB0_IO_066_mb1_FB1_TB2_IO_064,
    input wire        mb1_FA1_TB0_IO_067_mb1_FB1_TB2_IO_065,
    input wire        mb1_FA1_TB0_IO_068_mb1_FB1_TB2_IO_082,
    input wire        mb1_FA1_TB0_IO_069_mb1_FB1_TB2_IO_083,
    input wire        mb1_FA1_TB0_IO_070_mb1_FB1_TB2_IO_060,
    input wire        mb1_FA1_TB0_IO_071_mb1_FB1_TB2_IO_061,
    input wire        mb1_FA1_TB0_IO_072_mb1_FB1_TB2_IO_058,
    input wire        mb1_FA1_TB0_IO_073_mb1_FB1_TB2_IO_059,
    input wire        mb1_FA1_TB0_IO_074_mb1_FB1_TB2_IO_076,
    input wire        mb1_FA1_TB0_IO_075_mb1_FB1_TB2_IO_077,
    input wire        mb1_FA1_TB0_IO_076_mb1_FB1_TB2_IO_074,
    input wire        mb1_FA1_TB0_IO_077_mb1_FB1_TB2_IO_075,
    input wire        mb1_FA1_TB0_IO_078_mb1_FB1_TB2_IO_092,
    input wire        mb1_FA1_TB0_IO_079_mb1_FB1_TB2_IO_093,
    input wire        mb1_FA1_TB0_IO_080_mb1_FB1_TB2_IO_090,
    input wire        mb1_FA1_TB0_IO_081_mb1_FB1_TB2_IO_091,
    input wire        mb1_FA1_TB0_IO_082_mb1_FB1_TB2_IO_068,
    input wire        mb1_FA1_TB0_IO_083_mb1_FB1_TB2_IO_069,
    input wire        mb1_FA1_TB0_IO_084_mb1_FB1_TB2_IO_086,
    input wire        mb1_FA1_TB0_IO_085_mb1_FB1_TB2_IO_087,
    input wire        mb1_FA1_TB0_IO_086_mb1_FB1_TB2_IO_084,
    input wire        mb1_FA1_TB0_IO_087_mb1_FB1_TB2_IO_085,
    input wire        mb1_FA1_TB0_IO_088_mb1_FB1_TB2_IO_102,
    input wire        mb1_FA1_TB0_IO_089_mb1_FB1_TB2_IO_103,
    input wire        mb1_FA1_TB0_IO_090_mb1_FB1_TB2_IO_080,
    input wire        mb1_FA1_TB0_IO_091_mb1_FB1_TB2_IO_081,
    input wire        mb1_FA1_TB0_IO_092_mb1_FB1_TB2_IO_078,
    input wire        mb1_FA1_TB0_IO_093_mb1_FB1_TB2_IO_079,
    input wire        mb1_FA1_TB0_IO_094_mb1_FB1_TB2_IO_096,
    input wire        mb1_FA1_TB0_IO_095_mb1_FB1_TB2_IO_097,
    input wire        mb1_FA1_TB0_IO_096_mb1_FB1_TB2_IO_094,
    input wire        mb1_FA1_TB0_IO_097_mb1_FB1_TB2_IO_095,
    input wire        mb1_FA1_TB0_IO_098_mb1_FB1_TB2_IO_112,
    input wire        mb1_FA1_TB0_IO_099_mb1_FB1_TB2_IO_113,
    input wire        mb1_FA1_TB0_IO_100_mb1_FB1_TB2_IO_110,
    input wire        mb1_FA1_TB0_IO_101_mb1_FB1_TB2_IO_111,
    input wire        mb1_FA1_TB0_IO_102_mb1_FB1_TB2_IO_088,
    input wire        mb1_FA1_TB0_IO_103_mb1_FB1_TB2_IO_089,
    input wire        mb1_FA1_TB0_IO_104_mb1_FB1_TB2_IO_106,
    input wire        mb1_FA1_TB0_IO_105_mb1_FB1_TB2_IO_107,
    input wire        mb1_FA1_TB0_IO_106_mb1_FB1_TB2_IO_104,
    input wire        mb1_FA1_TB0_IO_107_mb1_FB1_TB2_IO_105,
    input wire        mb1_FA1_TB0_IO_108_mb1_FB1_TB2_IO_122,
    input wire        mb1_FA1_TB0_IO_109_mb1_FB1_TB2_IO_123,
    input wire        mb1_FA1_TB0_IO_110_mb1_FB1_TB2_IO_100,
    input wire        mb1_FA1_TB0_IO_111_mb1_FB1_TB2_IO_101,
    input wire        mb1_FA1_TB0_IO_112_mb1_FB1_TB2_IO_098,
    input wire        mb1_FA1_TB0_IO_113_mb1_FB1_TB2_IO_099,
    input wire        mb1_FA1_TB0_IO_114_mb1_FB1_TB2_IO_116,
    input wire        mb1_FA1_TB0_IO_115_mb1_FB1_TB2_IO_117,
    input wire        mb1_FA1_TB0_IO_116_mb1_FB1_TB2_IO_114,
    input wire        mb1_FA1_TB0_IO_117_mb1_FB1_TB2_IO_115,
    input wire        mb1_FA1_TB0_IO_118_mb1_FB1_TB2_IO_132,
    input wire        mb1_FA1_TB0_IO_119_mb1_FB1_TB2_IO_133,
    input wire        mb1_FA1_TB0_IO_120_mb1_FB1_TB2_IO_130,
    input wire        mb1_FA1_TB0_IO_121_mb1_FB1_TB2_IO_131,
    input wire        mb1_FA1_TB0_IO_122_mb1_FB1_TB2_IO_108,
    input wire        mb1_FA1_TB0_IO_123_mb1_FB1_TB2_IO_109,
    input wire        mb1_FA1_TB0_IO_124_mb1_FB1_TB2_IO_126,
    input wire        mb1_FA1_TB0_IO_125_mb1_FB1_TB2_IO_127,
    input wire        mb1_FA1_TB0_IO_126_mb1_FB1_TB2_IO_124,
    input wire        mb1_FA1_TB0_IO_127_mb1_FB1_TB2_IO_125,
    input wire        mb1_FA1_TB0_IO_130_mb1_FB1_TB2_IO_120,
    input wire        mb1_FA1_TB0_IO_131_mb1_FB1_TB2_IO_121,
    input wire        mb1_FA1_TB0_IO_132_mb1_FB1_TB2_IO_118,
    input wire        mb1_FA1_TB0_IO_133_mb1_FB1_TB2_IO_119,
    input wire        mb1_FA1_TB0_IO_134_mb1_FB1_TB2_IO_136,
    input wire        mb1_FA1_TB0_IO_136_mb1_FB1_TB2_IO_134,
    output wire        mb1_FB1_BA0_CLKIO_N_0_mb1_FA2_TB1_CLKIO_N_7,
    output wire        mb1_FB1_BA0_CLKIO_N_1_mb1_FA2_TB1_CLKIO_N_6,
    output wire        mb1_FB1_BA0_CLKIO_N_2_mb1_FA2_TB1_CLKIO_N_4,
    output wire        mb1_FB1_BA0_CLKIO_N_3_mb1_FA2_TB1_CLKIO_N_3,
    output wire        mb1_FB1_BA0_CLKIO_N_4_mb1_FA2_TB1_CLKIO_N_2,
    output wire        mb1_FB1_BA0_CLKIO_N_5_mb1_FA2_TB1_IO_010,
    output wire        mb1_FB1_BA0_CLKIO_N_6_mb1_FA2_TB1_CLKIO_N_1,
    output wire        mb1_FB1_BA0_CLKIO_N_7_mb1_FA2_TB1_CLKIO_N_0,
    output wire        mb1_FB1_BA0_CLKIO_P_0_mb1_FA2_TB1_CLKIO_P_7,
    output wire        mb1_FB1_BA0_CLKIO_P_1_mb1_FA2_TB1_CLKIO_P_6,
    output wire        mb1_FB1_BA0_CLKIO_P_2_mb1_FA2_TB1_CLKIO_P_4,
    output wire        mb1_FB1_BA0_CLKIO_P_3_mb1_FA2_TB1_CLKIO_P_3,
    output wire        mb1_FB1_BA0_CLKIO_P_4_mb1_FA2_TB1_CLKIO_P_2,
    output wire        mb1_FB1_BA0_CLKIO_P_5_mb1_FA2_TB1_IO_011,
    output wire        mb1_FB1_BA0_CLKIO_P_6_mb1_FA2_TB1_CLKIO_P_1,
    output wire        mb1_FB1_BA0_CLKIO_P_7_mb1_FA2_TB1_CLKIO_P_0,
    output wire        mb1_FB1_BA0_IO_004_mb1_FA2_TB1_IO_006,
    output wire        mb1_FB1_BA0_IO_005_mb1_FA2_TB1_IO_007,
    output wire        mb1_FB1_BA0_IO_006_mb1_FA2_TB1_IO_004,
    output wire        mb1_FB1_BA0_IO_007_mb1_FA2_TB1_IO_005,
    output wire        mb1_FB1_BA0_IO_008_mb1_FA2_TB1_IO_022,
    output wire        mb1_FB1_BA0_IO_009_mb1_FA2_TB1_IO_023,
    output wire        mb1_FB1_BA0_IO_010_mb1_FA2_TB1_CLKIO_N_5,
    output wire        mb1_FB1_BA0_IO_011_mb1_FA2_TB1_CLKIO_P_5,
    output wire        mb1_FB1_BA0_IO_012_mb1_FA2_TB1_IO_012,
    output wire        mb1_FB1_BA0_IO_013_mb1_FA2_TB1_IO_013,
    output wire        mb1_FB1_BA0_IO_014_mb1_FA2_TB1_IO_016,
    output wire        mb1_FB1_BA0_IO_015_mb1_FA2_TB1_IO_017,
    output wire        mb1_FB1_BA0_IO_016_mb1_FA2_TB1_IO_014,
    output wire        mb1_FB1_BA0_IO_017_mb1_FA2_TB1_IO_015,
    output wire        mb1_FB1_BA0_IO_018_mb1_FA2_TB1_IO_032,
    output wire        mb1_FB1_BA0_IO_019_mb1_FA2_TB1_IO_033,
    output wire        mb1_FB1_BA0_IO_020_mb1_FA2_TB1_IO_030,
    output wire        mb1_FB1_BA0_IO_021_mb1_FA2_TB1_IO_031,
    output wire        mb1_FB1_BA0_IO_022_mb1_FA2_TB1_IO_008,
    output wire        mb1_FB1_BA0_IO_023_mb1_FA2_TB1_IO_009,
    output wire        mb1_FB1_BA0_IO_024_mb1_FA2_TB1_IO_026,
    output wire        mb1_FB1_BA0_IO_025_mb1_FA2_TB1_IO_027,
    output wire        mb1_FB1_BA0_IO_026_mb1_FA2_TB1_IO_024,
    output wire        mb1_FB1_BA0_IO_027_mb1_FA2_TB1_IO_025,
    output wire        mb1_FB1_BA0_IO_028_mb1_FA2_TB1_IO_042,
    output wire        mb1_FB1_BA0_IO_029_mb1_FA2_TB1_IO_043,
    output wire        mb1_FB1_BA0_IO_030_mb1_FA2_TB1_IO_020,
    output wire        mb1_FB1_BA0_IO_031_mb1_FA2_TB1_IO_021,
    output wire        mb1_FB1_BA0_IO_032_mb1_FA2_TB1_IO_018,
    output wire        mb1_FB1_BA0_IO_033_mb1_FA2_TB1_IO_019,
    output wire        mb1_FB1_BA0_IO_034_mb1_FA2_TB1_IO_036,
    output wire        mb1_FB1_BA0_IO_035_mb1_FA2_TB1_IO_037,
    output wire        mb1_FB1_BA0_IO_036_mb1_FA2_TB1_IO_034,
    output wire        mb1_FB1_BA0_IO_037_mb1_FA2_TB1_IO_035,
    output wire        mb1_FB1_BA0_IO_038_mb1_FA2_TB1_IO_052,
    output wire        mb1_FB1_BA0_IO_039_mb1_FA2_TB1_IO_053,
    output wire        mb1_FB1_BA0_IO_040_mb1_FA2_TB1_IO_050,
    output wire        mb1_FB1_BA0_IO_041_mb1_FA2_TB1_IO_051,
    output wire        mb1_FB1_BA0_IO_042_mb1_FA2_TB1_IO_028,
    output wire        mb1_FB1_BA0_IO_043_mb1_FA2_TB1_IO_029,
    output wire        mb1_FB1_BA0_IO_044_mb1_FA2_TB1_IO_046,
    output wire        mb1_FB1_BA0_IO_045_mb1_FA2_TB1_IO_047,
    output wire        mb1_FB1_BA0_IO_046_mb1_FA2_TB1_IO_044,
    output wire        mb1_FB1_BA0_IO_047_mb1_FA2_TB1_IO_045,
    output wire        mb1_FB1_BA0_IO_048_mb1_FA2_TB1_IO_062,
    output wire        mb1_FB1_BA0_IO_049_mb1_FA2_TB1_IO_063,
    output wire        mb1_FB1_BA0_IO_050_mb1_FA2_TB1_IO_040,
    output wire        mb1_FB1_BA0_IO_051_mb1_FA2_TB1_IO_041,
    output wire        mb1_FB1_BA0_IO_052_mb1_FA2_TB1_IO_038,
    output wire        mb1_FB1_BA0_IO_053_mb1_FA2_TB1_IO_039,
    output wire        mb1_FB1_BA0_IO_054_mb1_FA2_TB1_IO_056,
    output wire        mb1_FB1_BA0_IO_055_mb1_FA2_TB1_IO_057,
    output wire        mb1_FB1_BA0_IO_056_mb1_FA2_TB1_IO_054,
    output wire        mb1_FB1_BA0_IO_057_mb1_FA2_TB1_IO_055,
    output wire        mb1_FB1_BA0_IO_058_mb1_FA2_TB1_IO_072,
    output wire        mb1_FB1_BA0_IO_059_mb1_FA2_TB1_IO_073,
    output wire        mb1_FB1_BA0_IO_060_mb1_FA2_TB1_IO_070,
    output wire        mb1_FB1_BA0_IO_061_mb1_FA2_TB1_IO_071,
    output wire        mb1_FB1_BA0_IO_062_mb1_FA2_TB1_IO_048,
    output wire        mb1_FB1_BA0_IO_063_mb1_FA2_TB1_IO_049,
    output wire        mb1_FB1_BA0_IO_064_mb1_FA2_TB1_IO_066,
    output wire        mb1_FB1_BA0_IO_065_mb1_FA2_TB1_IO_067,
    output wire        mb1_FB1_BA0_IO_066_mb1_FA2_TB1_IO_064,
    output wire        mb1_FB1_BA0_IO_067_mb1_FA2_TB1_IO_065,
    output wire        mb1_FB1_BA0_IO_068_mb1_FA2_TB1_IO_082,
    output wire        mb1_FB1_BA0_IO_069_mb1_FA2_TB1_IO_083,
    output wire        mb1_FB1_BA0_IO_070_mb1_FA2_TB1_IO_060,
    output wire        mb1_FB1_BA0_IO_071_mb1_FA2_TB1_IO_061,
    output wire        mb1_FB1_BA0_IO_072_mb1_FA2_TB1_IO_058,
    output wire        mb1_FB1_BA0_IO_073_mb1_FA2_TB1_IO_059,
    output wire        mb1_FB1_BA0_IO_074_mb1_FA2_TB1_IO_076,
    output wire        mb1_FB1_BA0_IO_075_mb1_FA2_TB1_IO_077,
    output wire        mb1_FB1_BA0_IO_076_mb1_FA2_TB1_IO_074,
    output wire        mb1_FB1_BA0_IO_077_mb1_FA2_TB1_IO_075,
    output wire        mb1_FB1_BA0_IO_078_mb1_FA2_TB1_IO_092,
    output wire        mb1_FB1_BA0_IO_079_mb1_FA2_TB1_IO_093,
    output wire        mb1_FB1_BA0_IO_080_mb1_FA2_TB1_IO_090,
    output wire        mb1_FB1_BA0_IO_081_mb1_FA2_TB1_IO_091,
    output wire        mb1_FB1_BA0_IO_082_mb1_FA2_TB1_IO_068,
    output wire        mb1_FB1_BA0_IO_083_mb1_FA2_TB1_IO_069,
    output wire        mb1_FB1_BA0_IO_084_mb1_FA2_TB1_IO_086,
    output wire        mb1_FB1_BA0_IO_085_mb1_FA2_TB1_IO_087,
    output wire        mb1_FB1_BA0_IO_086_mb1_FA2_TB1_IO_084,
    output wire        mb1_FB1_BA0_IO_087_mb1_FA2_TB1_IO_085,
    output wire        mb1_FB1_BA0_IO_088_mb1_FA2_TB1_IO_102,
    output wire        mb1_FB1_BA0_IO_089_mb1_FA2_TB1_IO_103,
    output wire        mb1_FB1_BA0_IO_090_mb1_FA2_TB1_IO_080,
    output wire        mb1_FB1_BA0_IO_091_mb1_FA2_TB1_IO_081,
    output wire        mb1_FB1_BA0_IO_092_mb1_FA2_TB1_IO_078,
    output wire        mb1_FB1_BA0_IO_093_mb1_FA2_TB1_IO_079,
    output wire        mb1_FB1_BA0_IO_094_mb1_FA2_TB1_IO_096,
    output wire        mb1_FB1_BA0_IO_095_mb1_FA2_TB1_IO_097,
    output wire        mb1_FB1_BA0_IO_096_mb1_FA2_TB1_IO_094,
    output wire        mb1_FB1_BA0_IO_097_mb1_FA2_TB1_IO_095,
    output wire        mb1_FB1_BA0_IO_098_mb1_FA2_TB1_IO_112,
    output wire        mb1_FB1_BA0_IO_099_mb1_FA2_TB1_IO_113,
    output wire        mb1_FB1_BA0_IO_100_mb1_FA2_TB1_IO_110,
    output wire        mb1_FB1_BA0_IO_101_mb1_FA2_TB1_IO_111,
    output wire        mb1_FB1_BA0_IO_102_mb1_FA2_TB1_IO_088,
    output wire        mb1_FB1_BA0_IO_103_mb1_FA2_TB1_IO_089,
    output wire        mb1_FB1_BA0_IO_104_mb1_FA2_TB1_IO_106,
    output wire        mb1_FB1_BA0_IO_105_mb1_FA2_TB1_IO_107,
    output wire        mb1_FB1_BA0_IO_106_mb1_FA2_TB1_IO_104,
    output wire        mb1_FB1_BA0_IO_107_mb1_FA2_TB1_IO_105,
    output wire        mb1_FB1_BA0_IO_108_mb1_FA2_TB1_IO_122,
    output wire        mb1_FB1_BA0_IO_109_mb1_FA2_TB1_IO_123,
    output wire        mb1_FB1_BA0_IO_110_mb1_FA2_TB1_IO_100,
    output wire        mb1_FB1_BA0_IO_111_mb1_FA2_TB1_IO_101,
    output wire        mb1_FB1_BA0_IO_112_mb1_FA2_TB1_IO_098,
    output wire        mb1_FB1_BA0_IO_113_mb1_FA2_TB1_IO_099,
    output wire        mb1_FB1_BA0_IO_114_mb1_FA2_TB1_IO_116,
    output wire        mb1_FB1_BA0_IO_115_mb1_FA2_TB1_IO_117,
    output wire        mb1_FB1_BA0_IO_116_mb1_FA2_TB1_IO_114,
    output wire        mb1_FB1_BA0_IO_117_mb1_FA2_TB1_IO_115,
    output wire        mb1_FB1_BA0_IO_118_mb1_FA2_TB1_IO_132,
    output wire        mb1_FB1_BA0_IO_119_mb1_FA2_TB1_IO_133,
    output wire        mb1_FB1_BA0_IO_120_mb1_FA2_TB1_IO_130,
    output wire        mb1_FB1_BA0_IO_121_mb1_FA2_TB1_IO_131,
    output wire        mb1_FB1_BA0_IO_122_mb1_FA2_TB1_IO_108,
    output wire        mb1_FB1_BA0_IO_123_mb1_FA2_TB1_IO_109,
    output wire        mb1_FB1_BA0_IO_124_mb1_FA2_TB1_IO_126,
    output wire        mb1_FB1_BA0_IO_125_mb1_FA2_TB1_IO_127,
    output wire        mb1_FB1_BA0_IO_126_mb1_FA2_TB1_IO_124,
    output wire        mb1_FB1_BA0_IO_127_mb1_FA2_TB1_IO_125,
    output wire        mb1_FB1_BA0_IO_130_mb1_FA2_TB1_IO_120,
    output wire        mb1_FB1_BA0_IO_131_mb1_FA2_TB1_IO_121,
    output wire        mb1_FB1_BA0_IO_132_mb1_FA2_TB1_IO_118,
    output wire        mb1_FB1_BA0_IO_133_mb1_FA2_TB1_IO_119,
    output wire        mb1_FB1_BA0_IO_134_mb1_FA2_TB1_IO_136,
    output wire        mb1_FB1_BA0_IO_136_mb1_FA2_TB1_IO_134,
    output wire        mb1_FB1_BA1_CLKIO_N_0_mb1_FA2_TB0_CLKIO_N_7,
    output wire        mb1_FB1_BA1_CLKIO_N_1_mb1_FA2_TB0_CLKIO_N_6,
    output wire        mb1_FB1_BA1_CLKIO_N_2_mb1_FA2_TB0_CLKIO_N_4,
    output wire        mb1_FB1_BA1_CLKIO_N_3_mb1_FA2_TB0_CLKIO_N_3,
    output wire        mb1_FB1_BA1_CLKIO_N_4_mb1_FA2_TB0_CLKIO_N_2,
    output wire        mb1_FB1_BA1_CLKIO_N_5_mb1_FA2_TB0_IO_010,
    output wire        mb1_FB1_BA1_CLKIO_N_6_mb1_FA2_TB0_CLKIO_N_1,
    output wire        mb1_FB1_BA1_CLKIO_N_7_mb1_FA2_TB0_CLKIO_N_0,
    output wire        mb1_FB1_BA1_CLKIO_P_0_mb1_FA2_TB0_CLKIO_P_7,
    output wire        mb1_FB1_BA1_CLKIO_P_1_mb1_FA2_TB0_CLKIO_P_6,
    output wire        mb1_FB1_BA1_CLKIO_P_2_mb1_FA2_TB0_CLKIO_P_4,
    output wire        mb1_FB1_BA1_CLKIO_P_3_mb1_FA2_TB0_CLKIO_P_3,
    output wire        mb1_FB1_BA1_CLKIO_P_4_mb1_FA2_TB0_CLKIO_P_2,
    output wire        mb1_FB1_BA1_CLKIO_P_5_mb1_FA2_TB0_IO_011,
    output wire        mb1_FB1_BA1_CLKIO_P_6_mb1_FA2_TB0_CLKIO_P_1,
    output wire        mb1_FB1_BA1_CLKIO_P_7_mb1_FA2_TB0_CLKIO_P_0,
    output wire        mb1_FB1_BA1_IO_004_mb1_FA2_TB0_IO_006,
    output wire        mb1_FB1_BA1_IO_005_mb1_FA2_TB0_IO_007,
    output wire        mb1_FB1_BA1_IO_006_mb1_FA2_TB0_IO_004,
    output wire        mb1_FB1_BA1_IO_007_mb1_FA2_TB0_IO_005,
    output wire        mb1_FB1_BA1_IO_008_mb1_FA2_TB0_IO_022,
    output wire        mb1_FB1_BA1_IO_009_mb1_FA2_TB0_IO_023,
    output wire        mb1_FB1_BA1_IO_010_mb1_FA2_TB0_CLKIO_N_5,
    output wire        mb1_FB1_BA1_IO_011_mb1_FA2_TB0_CLKIO_P_5,
    output wire        mb1_FB1_BA1_IO_012_mb1_FA2_TB0_IO_012,
    output wire        mb1_FB1_BA1_IO_013_mb1_FA2_TB0_IO_013,
    output wire        mb1_FB1_BA1_IO_014_mb1_FA2_TB0_IO_016,
    output wire        mb1_FB1_BA1_IO_015_mb1_FA2_TB0_IO_017,
    output wire        mb1_FB1_BA1_IO_016_mb1_FA2_TB0_IO_014,
    output wire        mb1_FB1_BA1_IO_017_mb1_FA2_TB0_IO_015,
    output wire        mb1_FB1_BA1_IO_018_mb1_FA2_TB0_IO_032,
    output wire        mb1_FB1_BA1_IO_019_mb1_FA2_TB0_IO_033,
    output wire        mb1_FB1_BA1_IO_020_mb1_FA2_TB0_IO_030,
    output wire        mb1_FB1_BA1_IO_021_mb1_FA2_TB0_IO_031,
    output wire        mb1_FB1_BA1_IO_022_mb1_FA2_TB0_IO_008,
    output wire        mb1_FB1_BA1_IO_023_mb1_FA2_TB0_IO_009,
    output wire        mb1_FB1_BA1_IO_024_mb1_FA2_TB0_IO_026,
    output wire        mb1_FB1_BA1_IO_025_mb1_FA2_TB0_IO_027,
    output wire        mb1_FB1_BA1_IO_026_mb1_FA2_TB0_IO_024,
    output wire        mb1_FB1_BA1_IO_027_mb1_FA2_TB0_IO_025,
    output wire        mb1_FB1_BA1_IO_028_mb1_FA2_TB0_IO_042,
    output wire        mb1_FB1_BA1_IO_029_mb1_FA2_TB0_IO_043,
    output wire        mb1_FB1_BA1_IO_030_mb1_FA2_TB0_IO_020,
    output wire        mb1_FB1_BA1_IO_031_mb1_FA2_TB0_IO_021,
    output wire        mb1_FB1_BA1_IO_032_mb1_FA2_TB0_IO_018,
    output wire        mb1_FB1_BA1_IO_033_mb1_FA2_TB0_IO_019,
    output wire        mb1_FB1_BA1_IO_034_mb1_FA2_TB0_IO_036,
    output wire        mb1_FB1_BA1_IO_035_mb1_FA2_TB0_IO_037,
    output wire        mb1_FB1_BA1_IO_036_mb1_FA2_TB0_IO_034,
    output wire        mb1_FB1_BA1_IO_037_mb1_FA2_TB0_IO_035,
    output wire        mb1_FB1_BA1_IO_038_mb1_FA2_TB0_IO_052,
    output wire        mb1_FB1_BA1_IO_039_mb1_FA2_TB0_IO_053,
    output wire        mb1_FB1_BA1_IO_040_mb1_FA2_TB0_IO_050,
    output wire        mb1_FB1_BA1_IO_041_mb1_FA2_TB0_IO_051,
    output wire        mb1_FB1_BA1_IO_042_mb1_FA2_TB0_IO_028,
    output wire        mb1_FB1_BA1_IO_043_mb1_FA2_TB0_IO_029,
    output wire        mb1_FB1_BA1_IO_044_mb1_FA2_TB0_IO_046,
    output wire        mb1_FB1_BA1_IO_045_mb1_FA2_TB0_IO_047,
    output wire        mb1_FB1_BA1_IO_046_mb1_FA2_TB0_IO_044,
    output wire        mb1_FB1_BA1_IO_047_mb1_FA2_TB0_IO_045,
    output wire        mb1_FB1_BA1_IO_048_mb1_FA2_TB0_IO_062,
    output wire        mb1_FB1_BA1_IO_049_mb1_FA2_TB0_IO_063,
    output wire        mb1_FB1_BA1_IO_050_mb1_FA2_TB0_IO_040,
    output wire        mb1_FB1_BA1_IO_051_mb1_FA2_TB0_IO_041,
    output wire        mb1_FB1_BA1_IO_052_mb1_FA2_TB0_IO_038,
    output wire        mb1_FB1_BA1_IO_053_mb1_FA2_TB0_IO_039,
    output wire        mb1_FB1_BA1_IO_054_mb1_FA2_TB0_IO_056,
    output wire        mb1_FB1_BA1_IO_055_mb1_FA2_TB0_IO_057,
    output wire        mb1_FB1_BA1_IO_056_mb1_FA2_TB0_IO_054,
    output wire        mb1_FB1_BA1_IO_057_mb1_FA2_TB0_IO_055,
    output wire        mb1_FB1_BA1_IO_058_mb1_FA2_TB0_IO_072,
    output wire        mb1_FB1_BA1_IO_059_mb1_FA2_TB0_IO_073,
    output wire        mb1_FB1_BA1_IO_060_mb1_FA2_TB0_IO_070,
    output wire        mb1_FB1_BA1_IO_061_mb1_FA2_TB0_IO_071,
    output wire        mb1_FB1_BA1_IO_062_mb1_FA2_TB0_IO_048,
    output wire        mb1_FB1_BA1_IO_063_mb1_FA2_TB0_IO_049,
    output wire        mb1_FB1_BA1_IO_064_mb1_FA2_TB0_IO_066,
    output wire        mb1_FB1_BA1_IO_065_mb1_FA2_TB0_IO_067,
    output wire        mb1_FB1_BA1_IO_066_mb1_FA2_TB0_IO_064,
    output wire        mb1_FB1_BA1_IO_067_mb1_FA2_TB0_IO_065,
    output wire        mb1_FB1_BA1_IO_068_mb1_FA2_TB0_IO_082,
    output wire        mb1_FB1_BA1_IO_069_mb1_FA2_TB0_IO_083,
    output wire        mb1_FB1_BA1_IO_070_mb1_FA2_TB0_IO_060,
    output wire        mb1_FB1_BA1_IO_071_mb1_FA2_TB0_IO_061,
    output wire        mb1_FB1_BA1_IO_072_mb1_FA2_TB0_IO_058,
    output wire        mb1_FB1_BA1_IO_073_mb1_FA2_TB0_IO_059,
    output wire        mb1_FB1_BA1_IO_074_mb1_FA2_TB0_IO_076,
    output wire        mb1_FB1_BA1_IO_075_mb1_FA2_TB0_IO_077,
    output wire        mb1_FB1_BA1_IO_076_mb1_FA2_TB0_IO_074,
    output wire        mb1_FB1_BA1_IO_077_mb1_FA2_TB0_IO_075,
    output wire        mb1_FB1_BA1_IO_078_mb1_FA2_TB0_IO_092,
    output wire        mb1_FB1_BA1_IO_079_mb1_FA2_TB0_IO_093,
    output wire        mb1_FB1_BA1_IO_080_mb1_FA2_TB0_IO_090,
    output wire        mb1_FB1_BA1_IO_081_mb1_FA2_TB0_IO_091,
    output wire        mb1_FB1_BA1_IO_082_mb1_FA2_TB0_IO_068,
    output wire        mb1_FB1_BA1_IO_083_mb1_FA2_TB0_IO_069,
    output wire        mb1_FB1_BA1_IO_084_mb1_FA2_TB0_IO_086,
    output wire        mb1_FB1_BA1_IO_085_mb1_FA2_TB0_IO_087,
    output wire        mb1_FB1_BA1_IO_086_mb1_FA2_TB0_IO_084,
    output wire        mb1_FB1_BA1_IO_087_mb1_FA2_TB0_IO_085,
    output wire        mb1_FB1_BA1_IO_088_mb1_FA2_TB0_IO_102,
    output wire        mb1_FB1_BA1_IO_089_mb1_FA2_TB0_IO_103,
    output wire        mb1_FB1_BA1_IO_090_mb1_FA2_TB0_IO_080,
    output wire        mb1_FB1_BA1_IO_091_mb1_FA2_TB0_IO_081,
    output wire        mb1_FB1_BA1_IO_092_mb1_FA2_TB0_IO_078,
    output wire        mb1_FB1_BA1_IO_093_mb1_FA2_TB0_IO_079,
    output wire        mb1_FB1_BA1_IO_094_mb1_FA2_TB0_IO_096,
    output wire        mb1_FB1_BA1_IO_095_mb1_FA2_TB0_IO_097,
    output wire        mb1_FB1_BA1_IO_096_mb1_FA2_TB0_IO_094,
    output wire        mb1_FB1_BA1_IO_097_mb1_FA2_TB0_IO_095,
    output wire        mb1_FB1_BA1_IO_098_mb1_FA2_TB0_IO_112,
    output wire        mb1_FB1_BA1_IO_099_mb1_FA2_TB0_IO_113,
    output wire        mb1_FB1_BA1_IO_100_mb1_FA2_TB0_IO_110,
    output wire        mb1_FB1_BA1_IO_101_mb1_FA2_TB0_IO_111,
    output wire        mb1_FB1_BA1_IO_102_mb1_FA2_TB0_IO_088,
    output wire        mb1_FB1_BA1_IO_103_mb1_FA2_TB0_IO_089,
    output wire        mb1_FB1_BA1_IO_104_mb1_FA2_TB0_IO_106,
    output wire        mb1_FB1_BA1_IO_105_mb1_FA2_TB0_IO_107,
    output wire        mb1_FB1_BA1_IO_106_mb1_FA2_TB0_IO_104,
    output wire        mb1_FB1_BA1_IO_107_mb1_FA2_TB0_IO_105,
    output wire        mb1_FB1_BA1_IO_108_mb1_FA2_TB0_IO_122,
    output wire        mb1_FB1_BA1_IO_109_mb1_FA2_TB0_IO_123,
    output wire        mb1_FB1_BA1_IO_110_mb1_FA2_TB0_IO_100,
    output wire        mb1_FB1_BA1_IO_111_mb1_FA2_TB0_IO_101,
    output wire        mb1_FB1_BA1_IO_112_mb1_FA2_TB0_IO_098,
    output wire        mb1_FB1_BA1_IO_113_mb1_FA2_TB0_IO_099,
    output wire        mb1_FB1_BA1_IO_114_mb1_FA2_TB0_IO_116,
    output wire        mb1_FB1_BA1_IO_115_mb1_FA2_TB0_IO_117,
    output wire        mb1_FB1_BA1_IO_116_mb1_FA2_TB0_IO_114,
    output wire        mb1_FB1_BA1_IO_117_mb1_FA2_TB0_IO_115,
    output wire        mb1_FB1_BA1_IO_118_mb1_FA2_TB0_IO_132,
    output wire        mb1_FB1_BA1_IO_119_mb1_FA2_TB0_IO_133,
    output wire        mb1_FB1_BA1_IO_120_mb1_FA2_TB0_IO_130,
    output wire        mb1_FB1_BA1_IO_121_mb1_FA2_TB0_IO_131,
    output wire        mb1_FB1_BA1_IO_122_mb1_FA2_TB0_IO_108,
    output wire        mb1_FB1_BA1_IO_123_mb1_FA2_TB0_IO_109,
    output wire        mb1_FB1_BA1_IO_124_mb1_FA2_TB0_IO_126,
    output wire        mb1_FB1_BA1_IO_125_mb1_FA2_TB0_IO_127,
    output wire        mb1_FB1_BA1_IO_126_mb1_FA2_TB0_IO_124,
    output wire        mb1_FB1_BA1_IO_127_mb1_FA2_TB0_IO_125,
    output wire        mb1_FB1_BA1_IO_130_mb1_FA2_TB0_IO_120,
    output wire        mb1_FB1_BA1_IO_131_mb1_FA2_TB0_IO_121,
    output wire        mb1_FB1_BA1_IO_132_mb1_FA2_TB0_IO_118,
    output wire        mb1_FB1_BA1_IO_133_mb1_FA2_TB0_IO_119,
    output wire        mb1_FB1_BA1_IO_134_mb1_FA2_TB0_IO_136,
    output wire        mb1_FB1_BA1_IO_136_mb1_FA2_TB0_IO_134,
    input wire        mb1_FA1_BA0_CLKIO_N_0_mb1_FB1_BA2_CLKIO_N_7,
    input wire        mb1_FA1_BA0_CLKIO_N_1_mb1_FB1_BA2_CLKIO_N_6,
    input wire        mb1_FA1_BA0_CLKIO_N_2_mb1_FB1_BA2_CLKIO_N_4,
    input wire        mb1_FA1_BA0_CLKIO_N_3_mb1_FB1_BA2_CLKIO_N_3,
    input wire        mb1_FA1_BA0_CLKIO_N_4_mb1_FB1_BA2_CLKIO_N_2,
    input wire        mb1_FA1_BA0_CLKIO_N_5_mb1_FB1_BA2_IO_010,
    input wire        mb1_FA1_BA0_CLKIO_N_6_mb1_FB1_BA2_CLKIO_N_1,
    input wire        mb1_FA1_BA0_CLKIO_N_7_mb1_FB1_BA2_CLKIO_N_0,
    input wire        mb1_FA1_BA0_CLKIO_P_0_mb1_FB1_BA2_CLKIO_P_7,
    input wire        mb1_FA1_BA0_CLKIO_P_1_mb1_FB1_BA2_CLKIO_P_6,
    input wire        mb1_FA1_BA0_CLKIO_P_2_mb1_FB1_BA2_CLKIO_P_4,
    input wire        mb1_FA1_BA0_CLKIO_P_3_mb1_FB1_BA2_CLKIO_P_3,
    input wire        mb1_FA1_BA0_CLKIO_P_4_mb1_FB1_BA2_CLKIO_P_2,
    input wire        mb1_FA1_BA0_CLKIO_P_5_mb1_FB1_BA2_IO_011,
    input wire        mb1_FA1_BA0_CLKIO_P_6_mb1_FB1_BA2_CLKIO_P_1,
    input wire        mb1_FA1_BA0_CLKIO_P_7_mb1_FB1_BA2_CLKIO_P_0,
    input wire        mb1_FA1_BA0_IO_004_mb1_FB1_BA2_IO_006,
    input wire        mb1_FA1_BA0_IO_005_mb1_FB1_BA2_IO_007,
    input wire        mb1_FA1_BA0_IO_006_mb1_FB1_BA2_IO_004,
    input wire        mb1_FA1_BA0_IO_007_mb1_FB1_BA2_IO_005,
    input wire        mb1_FA1_BA0_IO_008_mb1_FB1_BA2_IO_022,
    input wire        mb1_FA1_BA0_IO_009_mb1_FB1_BA2_IO_023,
    input wire        mb1_FA1_BA0_IO_010_mb1_FB1_BA2_CLKIO_N_5,
    input wire        mb1_FA1_BA0_IO_011_mb1_FB1_BA2_CLKIO_P_5,
    input wire        mb1_FA1_BA0_IO_012_mb1_FB1_BA2_IO_012,
    input wire        mb1_FA1_BA0_IO_013_mb1_FB1_BA2_IO_013,
    input wire        mb1_FA1_BA0_IO_014_mb1_FB1_BA2_IO_016,
    input wire        mb1_FA1_BA0_IO_015_mb1_FB1_BA2_IO_017,
    input wire        mb1_FA1_BA0_IO_016_mb1_FB1_BA2_IO_014,
    input wire        mb1_FA1_BA0_IO_017_mb1_FB1_BA2_IO_015,
    input wire        mb1_FA1_BA0_IO_018_mb1_FB1_BA2_IO_032,
    input wire        mb1_FA1_BA0_IO_019_mb1_FB1_BA2_IO_033,
    input wire        mb1_FA1_BA0_IO_020_mb1_FB1_BA2_IO_030,
    input wire        mb1_FA1_BA0_IO_021_mb1_FB1_BA2_IO_031,
    input wire        mb1_FA1_BA0_IO_022_mb1_FB1_BA2_IO_008,
    input wire        mb1_FA1_BA0_IO_023_mb1_FB1_BA2_IO_009,
    input wire        mb1_FA1_BA0_IO_024_mb1_FB1_BA2_IO_026,
    input wire        mb1_FA1_BA0_IO_025_mb1_FB1_BA2_IO_027,
    input wire        mb1_FA1_BA0_IO_026_mb1_FB1_BA2_IO_024,
    input wire        mb1_FA1_BA0_IO_027_mb1_FB1_BA2_IO_025,
    input wire        mb1_FA1_BA0_IO_028_mb1_FB1_BA2_IO_042,
    input wire        mb1_FA1_BA0_IO_029_mb1_FB1_BA2_IO_043,
    input wire        mb1_FA1_BA0_IO_030_mb1_FB1_BA2_IO_020,
    input wire        mb1_FA1_BA0_IO_031_mb1_FB1_BA2_IO_021,
    input wire        mb1_FA1_BA0_IO_032_mb1_FB1_BA2_IO_018,
    input wire        mb1_FA1_BA0_IO_033_mb1_FB1_BA2_IO_019,
    input wire        mb1_FA1_BA0_IO_034_mb1_FB1_BA2_IO_036,
    input wire        mb1_FA1_BA0_IO_035_mb1_FB1_BA2_IO_037,
    input wire        mb1_FA1_BA0_IO_036_mb1_FB1_BA2_IO_034,
    input wire        mb1_FA1_BA0_IO_037_mb1_FB1_BA2_IO_035,
    input wire        mb1_FA1_BA0_IO_038_mb1_FB1_BA2_IO_052,
    input wire        mb1_FA1_BA0_IO_039_mb1_FB1_BA2_IO_053,
    input wire        mb1_FA1_BA0_IO_040_mb1_FB1_BA2_IO_050,
    input wire        mb1_FA1_BA0_IO_041_mb1_FB1_BA2_IO_051,
    input wire        mb1_FA1_BA0_IO_042_mb1_FB1_BA2_IO_028,
    input wire        mb1_FA1_BA0_IO_043_mb1_FB1_BA2_IO_029,
    input wire        mb1_FA1_BA0_IO_044_mb1_FB1_BA2_IO_046,
    input wire        mb1_FA1_BA0_IO_045_mb1_FB1_BA2_IO_047,
    input wire        mb1_FA1_BA0_IO_046_mb1_FB1_BA2_IO_044,
    input wire        mb1_FA1_BA0_IO_047_mb1_FB1_BA2_IO_045,
    input wire        mb1_FA1_BA0_IO_048_mb1_FB1_BA2_IO_062,
    input wire        mb1_FA1_BA0_IO_049_mb1_FB1_BA2_IO_063,
    input wire        mb1_FA1_BA0_IO_050_mb1_FB1_BA2_IO_040,
    input wire        mb1_FA1_BA0_IO_051_mb1_FB1_BA2_IO_041,
    input wire        mb1_FA1_BA0_IO_052_mb1_FB1_BA2_IO_038,
    input wire        mb1_FA1_BA0_IO_053_mb1_FB1_BA2_IO_039,
    input wire        mb1_FA1_BA0_IO_054_mb1_FB1_BA2_IO_056,
    input wire        mb1_FA1_BA0_IO_055_mb1_FB1_BA2_IO_057,
    input wire        mb1_FA1_BA0_IO_056_mb1_FB1_BA2_IO_054,
    input wire        mb1_FA1_BA0_IO_057_mb1_FB1_BA2_IO_055,
    input wire        mb1_FA1_BA0_IO_058_mb1_FB1_BA2_IO_072,
    input wire        mb1_FA1_BA0_IO_059_mb1_FB1_BA2_IO_073,
    input wire        mb1_FA1_BA0_IO_060_mb1_FB1_BA2_IO_070,
    input wire        mb1_FA1_BA0_IO_061_mb1_FB1_BA2_IO_071,
    input wire        mb1_FA1_BA0_IO_062_mb1_FB1_BA2_IO_048,
    input wire        mb1_FA1_BA0_IO_063_mb1_FB1_BA2_IO_049,
    input wire        mb1_FA1_BA0_IO_064_mb1_FB1_BA2_IO_066,
    input wire        mb1_FA1_BA0_IO_065_mb1_FB1_BA2_IO_067,
    input wire        mb1_FA1_BA0_IO_066_mb1_FB1_BA2_IO_064,
    input wire        mb1_FA1_BA0_IO_067_mb1_FB1_BA2_IO_065,
    input wire        mb1_FA1_BA0_IO_068_mb1_FB1_BA2_IO_082,
    input wire        mb1_FA1_BA0_IO_069_mb1_FB1_BA2_IO_083,
    input wire        mb1_FA1_BA0_IO_070_mb1_FB1_BA2_IO_060,
    input wire        mb1_FA1_BA0_IO_071_mb1_FB1_BA2_IO_061,
    input wire        mb1_FA1_BA0_IO_072_mb1_FB1_BA2_IO_058,
    input wire        mb1_FA1_BA0_IO_073_mb1_FB1_BA2_IO_059,
    input wire        mb1_FA1_BA0_IO_074_mb1_FB1_BA2_IO_076,
    input wire        mb1_FA1_BA0_IO_075_mb1_FB1_BA2_IO_077,
    input wire        mb1_FA1_BA0_IO_076_mb1_FB1_BA2_IO_074,
    input wire        mb1_FA1_BA0_IO_077_mb1_FB1_BA2_IO_075,
    input wire        mb1_FA1_BA0_IO_078_mb1_FB1_BA2_IO_092,
    input wire        mb1_FA1_BA0_IO_079_mb1_FB1_BA2_IO_093,
    input wire        mb1_FA1_BA0_IO_080_mb1_FB1_BA2_IO_090,
    input wire        mb1_FA1_BA0_IO_081_mb1_FB1_BA2_IO_091,
    input wire        mb1_FA1_BA0_IO_082_mb1_FB1_BA2_IO_068,
    input wire        mb1_FA1_BA0_IO_083_mb1_FB1_BA2_IO_069,
    input wire        mb1_FA1_BA0_IO_084_mb1_FB1_BA2_IO_086,
    input wire        mb1_FA1_BA0_IO_085_mb1_FB1_BA2_IO_087,
    input wire        mb1_FA1_BA0_IO_086_mb1_FB1_BA2_IO_084,
    input wire        mb1_FA1_BA0_IO_087_mb1_FB1_BA2_IO_085,
    input wire        mb1_FA1_BA0_IO_088_mb1_FB1_BA2_IO_102,
    input wire        mb1_FA1_BA0_IO_089_mb1_FB1_BA2_IO_103,
    input wire        mb1_FA1_BA0_IO_090_mb1_FB1_BA2_IO_080,
    input wire        mb1_FA1_BA0_IO_091_mb1_FB1_BA2_IO_081,
    input wire        mb1_FA1_BA0_IO_092_mb1_FB1_BA2_IO_078,
    input wire        mb1_FA1_BA0_IO_093_mb1_FB1_BA2_IO_079,
    input wire        mb1_FA1_BA0_IO_094_mb1_FB1_BA2_IO_096,
    input wire        mb1_FA1_BA0_IO_095_mb1_FB1_BA2_IO_097,
    input wire        mb1_FA1_BA0_IO_096_mb1_FB1_BA2_IO_094,
    input wire        mb1_FA1_BA0_IO_097_mb1_FB1_BA2_IO_095,
    input wire        mb1_FA1_BA0_IO_098_mb1_FB1_BA2_IO_112,
    input wire        mb1_FA1_BA0_IO_099_mb1_FB1_BA2_IO_113,
    input wire        mb1_FA1_BA0_IO_100_mb1_FB1_BA2_IO_110,
    input wire        mb1_FA1_BA0_IO_101_mb1_FB1_BA2_IO_111,
    input wire        mb1_FA1_BA0_IO_102_mb1_FB1_BA2_IO_088,
    input wire        mb1_FA1_BA0_IO_103_mb1_FB1_BA2_IO_089,
    input wire        mb1_FA1_BA0_IO_104_mb1_FB1_BA2_IO_106,
    input wire        mb1_FA1_BA0_IO_105_mb1_FB1_BA2_IO_107,
    input wire        mb1_FA1_BA0_IO_106_mb1_FB1_BA2_IO_104,
    input wire        mb1_FA1_BA0_IO_107_mb1_FB1_BA2_IO_105,
    input wire        mb1_FA1_BA0_IO_108_mb1_FB1_BA2_IO_122,
    input wire        mb1_FA1_BA0_IO_109_mb1_FB1_BA2_IO_123,
    input wire        mb1_FA1_BA0_IO_110_mb1_FB1_BA2_IO_100,
    input wire        mb1_FA1_BA0_IO_111_mb1_FB1_BA2_IO_101,
    input wire        mb1_FA1_BA0_IO_112_mb1_FB1_BA2_IO_098,
    input wire        mb1_FA1_BA0_IO_113_mb1_FB1_BA2_IO_099,
    input wire        mb1_FA1_BA0_IO_114_mb1_FB1_BA2_IO_116,
    input wire        mb1_FA1_BA0_IO_115_mb1_FB1_BA2_IO_117,
    input wire        mb1_FA1_BA0_IO_116_mb1_FB1_BA2_IO_114,
    input wire        mb1_FA1_BA0_IO_117_mb1_FB1_BA2_IO_115,
    input wire        mb1_FA1_BA0_IO_118_mb1_FB1_BA2_IO_132,
    input wire        mb1_FA1_BA0_IO_119_mb1_FB1_BA2_IO_133,
    input wire        mb1_FA1_BA0_IO_120_mb1_FB1_BA2_IO_130,
    input wire        mb1_FA1_BA0_IO_121_mb1_FB1_BA2_IO_131,
    input wire        mb1_FA1_BA0_IO_122_mb1_FB1_BA2_IO_108,
    input wire        mb1_FA1_BA0_IO_123_mb1_FB1_BA2_IO_109,
    input wire        mb1_FA1_BA0_IO_124_mb1_FB1_BA2_IO_126,
    input wire        mb1_FA1_BA0_IO_125_mb1_FB1_BA2_IO_127,
    input wire        mb1_FA1_BA0_IO_126_mb1_FB1_BA2_IO_124,
    input wire        mb1_FA1_BA0_IO_127_mb1_FB1_BA2_IO_125,
    input wire        mb1_FA1_BA0_IO_130_mb1_FB1_BA2_IO_120,
    input wire        mb1_FA1_BA0_IO_131_mb1_FB1_BA2_IO_121,
    input wire        mb1_FA1_BA0_IO_132_mb1_FB1_BA2_IO_118,
    input wire        mb1_FA1_BA0_IO_133_mb1_FB1_BA2_IO_119,
    input wire        mb1_FA1_BA0_IO_134_mb1_FB1_BA2_IO_136,
    input wire        mb1_FA1_BA0_IO_136_mb1_FB1_BA2_IO_134,
    input wire        mb1_FA1_BA2_CLKIO_N_0_mb1_FB1_BB0_CLKIO_N_7,
    input wire        mb1_FA1_BA2_CLKIO_N_1_mb1_FB1_BB0_CLKIO_N_6,
    input wire        mb1_FA1_BA2_CLKIO_N_2_mb1_FB1_BB0_CLKIO_N_4,
    input wire        mb1_FA1_BA2_CLKIO_N_3_mb1_FB1_BB0_CLKIO_N_3,
    input wire        mb1_FA1_BA2_CLKIO_N_4_mb1_FB1_BB0_CLKIO_N_2,
    input wire        mb1_FA1_BA2_CLKIO_N_5_mb1_FB1_BB0_IO_010,
    input wire        mb1_FA1_BA2_CLKIO_N_6_mb1_FB1_BB0_CLKIO_N_1,
    input wire        mb1_FA1_BA2_CLKIO_N_7_mb1_FB1_BB0_CLKIO_N_0,
    input wire        mb1_FA1_BA2_CLKIO_P_0_mb1_FB1_BB0_CLKIO_P_7,
    input wire        mb1_FA1_BA2_CLKIO_P_1_mb1_FB1_BB0_CLKIO_P_6,
    input wire        mb1_FA1_BA2_CLKIO_P_2_mb1_FB1_BB0_CLKIO_P_4,
    input wire        mb1_FA1_BA2_CLKIO_P_3_mb1_FB1_BB0_CLKIO_P_3,
    input wire        mb1_FA1_BA2_CLKIO_P_4_mb1_FB1_BB0_CLKIO_P_2,
    input wire        mb1_FA1_BA2_CLKIO_P_5_mb1_FB1_BB0_IO_011,
    input wire        mb1_FA1_BA2_CLKIO_P_6_mb1_FB1_BB0_CLKIO_P_1,
    input wire        mb1_FA1_BA2_CLKIO_P_7_mb1_FB1_BB0_CLKIO_P_0,
    input wire        mb1_FA1_BA2_IO_004_mb1_FB1_BB0_IO_006,
    input wire        mb1_FA1_BA2_IO_005_mb1_FB1_BB0_IO_007,
    input wire        mb1_FA1_BA2_IO_006_mb1_FB1_BB0_IO_004,
    input wire        mb1_FA1_BA2_IO_007_mb1_FB1_BB0_IO_005,
    input wire        mb1_FA1_BA2_IO_008_mb1_FB1_BB0_IO_022,
    input wire        mb1_FA1_BA2_IO_009_mb1_FB1_BB0_IO_023,
    input wire        mb1_FA1_BA2_IO_010_mb1_FB1_BB0_CLKIO_N_5,
    input wire        mb1_FA1_BA2_IO_011_mb1_FB1_BB0_CLKIO_P_5,
    input wire        mb1_FA1_BA2_IO_012_mb1_FB1_BB0_IO_012,
    input wire        mb1_FA1_BA2_IO_013_mb1_FB1_BB0_IO_013,
    input wire        mb1_FA1_BA2_IO_014_mb1_FB1_BB0_IO_016,
    input wire        mb1_FA1_BA2_IO_015_mb1_FB1_BB0_IO_017,
    input wire        mb1_FA1_BA2_IO_016_mb1_FB1_BB0_IO_014,
    input wire        mb1_FA1_BA2_IO_017_mb1_FB1_BB0_IO_015,
    input wire        mb1_FA1_BA2_IO_018_mb1_FB1_BB0_IO_032,
    input wire        mb1_FA1_BA2_IO_019_mb1_FB1_BB0_IO_033,
    input wire        mb1_FA1_BA2_IO_020_mb1_FB1_BB0_IO_030,
    input wire        mb1_FA1_BA2_IO_021_mb1_FB1_BB0_IO_031,
    input wire        mb1_FA1_BA2_IO_022_mb1_FB1_BB0_IO_008,
    input wire        mb1_FA1_BA2_IO_023_mb1_FB1_BB0_IO_009,
    input wire        mb1_FA1_BA2_IO_024_mb1_FB1_BB0_IO_026,
    input wire        mb1_FA1_BA2_IO_025_mb1_FB1_BB0_IO_027,
    input wire        mb1_FA1_BA2_IO_026_mb1_FB1_BB0_IO_024,
    input wire        mb1_FA1_BA2_IO_027_mb1_FB1_BB0_IO_025,
    input wire        mb1_FA1_BA2_IO_028_mb1_FB1_BB0_IO_042,
    input wire        mb1_FA1_BA2_IO_029_mb1_FB1_BB0_IO_043,
    input wire        mb1_FA1_BA2_IO_030_mb1_FB1_BB0_IO_020,
    input wire        mb1_FA1_BA2_IO_031_mb1_FB1_BB0_IO_021,
    input wire        mb1_FA1_BA2_IO_032_mb1_FB1_BB0_IO_018,
    input wire        mb1_FA1_BA2_IO_033_mb1_FB1_BB0_IO_019,
    input wire        mb1_FA1_BA2_IO_034_mb1_FB1_BB0_IO_036,
    input wire        mb1_FA1_BA2_IO_035_mb1_FB1_BB0_IO_037,
    input wire        mb1_FA1_BA2_IO_036_mb1_FB1_BB0_IO_034,
    input wire        mb1_FA1_BA2_IO_037_mb1_FB1_BB0_IO_035,
    input wire        mb1_FA1_BA2_IO_038_mb1_FB1_BB0_IO_052,
    input wire        mb1_FA1_BA2_IO_039_mb1_FB1_BB0_IO_053,
    input wire        mb1_FA1_BA2_IO_040_mb1_FB1_BB0_IO_050,
    input wire        mb1_FA1_BA2_IO_041_mb1_FB1_BB0_IO_051,
    input wire        mb1_FA1_BA2_IO_042_mb1_FB1_BB0_IO_028,
    input wire        mb1_FA1_BA2_IO_043_mb1_FB1_BB0_IO_029,
    input wire        mb1_FA1_BA2_IO_044_mb1_FB1_BB0_IO_046,
    input wire        mb1_FA1_BA2_IO_045_mb1_FB1_BB0_IO_047,
    input wire        mb1_FA1_BA2_IO_046_mb1_FB1_BB0_IO_044,
    input wire        mb1_FA1_BA2_IO_047_mb1_FB1_BB0_IO_045,
    input wire        mb1_FA1_BA2_IO_048_mb1_FB1_BB0_IO_062,
    input wire        mb1_FA1_BA2_IO_049_mb1_FB1_BB0_IO_063,
    input wire        mb1_FA1_BA2_IO_050_mb1_FB1_BB0_IO_040,
    input wire        mb1_FA1_BA2_IO_051_mb1_FB1_BB0_IO_041,
    input wire        mb1_FA1_BA2_IO_052_mb1_FB1_BB0_IO_038,
    input wire        mb1_FA1_BA2_IO_053_mb1_FB1_BB0_IO_039,
    input wire        mb1_FA1_BA2_IO_054_mb1_FB1_BB0_IO_056,
    input wire        mb1_FA1_BA2_IO_055_mb1_FB1_BB0_IO_057,
    input wire        mb1_FA1_BA2_IO_056_mb1_FB1_BB0_IO_054,
    input wire        mb1_FA1_BA2_IO_057_mb1_FB1_BB0_IO_055,
    input wire        mb1_FA1_BA2_IO_058_mb1_FB1_BB0_IO_072,
    input wire        mb1_FA1_BA2_IO_059_mb1_FB1_BB0_IO_073,
    input wire        mb1_FA1_BA2_IO_060_mb1_FB1_BB0_IO_070,
    input wire        mb1_FA1_BA2_IO_061_mb1_FB1_BB0_IO_071,
    input wire        mb1_FA1_BA2_IO_062_mb1_FB1_BB0_IO_048,
    input wire        mb1_FA1_BA2_IO_063_mb1_FB1_BB0_IO_049,
    input wire        mb1_FA1_BA2_IO_064_mb1_FB1_BB0_IO_066,
    input wire        mb1_FA1_BA2_IO_065_mb1_FB1_BB0_IO_067,
    input wire        mb1_FA1_BA2_IO_066_mb1_FB1_BB0_IO_064,
    input wire        mb1_FA1_BA2_IO_067_mb1_FB1_BB0_IO_065,
    input wire        mb1_FA1_BA2_IO_068_mb1_FB1_BB0_IO_082,
    input wire        mb1_FA1_BA2_IO_069_mb1_FB1_BB0_IO_083,
    input wire        mb1_FA1_BA2_IO_070_mb1_FB1_BB0_IO_060,
    input wire        mb1_FA1_BA2_IO_071_mb1_FB1_BB0_IO_061,
    input wire        mb1_FA1_BA2_IO_072_mb1_FB1_BB0_IO_058,
    input wire        mb1_FA1_BA2_IO_073_mb1_FB1_BB0_IO_059,
    input wire        mb1_FA1_BA2_IO_074_mb1_FB1_BB0_IO_076,
    input wire        mb1_FA1_BA2_IO_075_mb1_FB1_BB0_IO_077,
    input wire        mb1_FA1_BA2_IO_076_mb1_FB1_BB0_IO_074,
    input wire        mb1_FA1_BA2_IO_077_mb1_FB1_BB0_IO_075,
    input wire        mb1_FA1_BA2_IO_078_mb1_FB1_BB0_IO_092,
    input wire        mb1_FA1_BA2_IO_079_mb1_FB1_BB0_IO_093,
    input wire        mb1_FA1_BA2_IO_080_mb1_FB1_BB0_IO_090,
    input wire        mb1_FA1_BA2_IO_081_mb1_FB1_BB0_IO_091,
    input wire        mb1_FA1_BA2_IO_082_mb1_FB1_BB0_IO_068,
    input wire        mb1_FA1_BA2_IO_083_mb1_FB1_BB0_IO_069,
    input wire        mb1_FA1_BA2_IO_084_mb1_FB1_BB0_IO_086,
    input wire        mb1_FA1_BA2_IO_085_mb1_FB1_BB0_IO_087,
    input wire        mb1_FA1_BA2_IO_086_mb1_FB1_BB0_IO_084,
    input wire        mb1_FA1_BA2_IO_087_mb1_FB1_BB0_IO_085,
    input wire        mb1_FA1_BA2_IO_088_mb1_FB1_BB0_IO_102,
    input wire        mb1_FA1_BA2_IO_089_mb1_FB1_BB0_IO_103,
    input wire        mb1_FA1_BA2_IO_090_mb1_FB1_BB0_IO_080,
    input wire        mb1_FA1_BA2_IO_091_mb1_FB1_BB0_IO_081,
    input wire        mb1_FA1_BA2_IO_092_mb1_FB1_BB0_IO_078,
    input wire        mb1_FA1_BA2_IO_093_mb1_FB1_BB0_IO_079,
    input wire        mb1_FA1_BA2_IO_094_mb1_FB1_BB0_IO_096,
    input wire        mb1_FA1_BA2_IO_095_mb1_FB1_BB0_IO_097,
    input wire        mb1_FA1_BA2_IO_096_mb1_FB1_BB0_IO_094,
    input wire        mb1_FA1_BA2_IO_097_mb1_FB1_BB0_IO_095,
    input wire        mb1_FA1_BA2_IO_098_mb1_FB1_BB0_IO_112,
    input wire        mb1_FA1_BA2_IO_099_mb1_FB1_BB0_IO_113,
    input wire        mb1_FA1_BA2_IO_100_mb1_FB1_BB0_IO_110,
    input wire        mb1_FA1_BA2_IO_101_mb1_FB1_BB0_IO_111,
    input wire        mb1_FA1_BA2_IO_102_mb1_FB1_BB0_IO_088,
    input wire        mb1_FA1_BA2_IO_103_mb1_FB1_BB0_IO_089,
    input wire        mb1_FA1_BA2_IO_104_mb1_FB1_BB0_IO_106,
    input wire        mb1_FA1_BA2_IO_105_mb1_FB1_BB0_IO_107,
    input wire        mb1_FA1_BA2_IO_106_mb1_FB1_BB0_IO_104,
    input wire        mb1_FA1_BA2_IO_107_mb1_FB1_BB0_IO_105,
    input wire        mb1_FA1_BA2_IO_108_mb1_FB1_BB0_IO_122,
    input wire        mb1_FA1_BA2_IO_109_mb1_FB1_BB0_IO_123,
    input wire        mb1_FA1_BA2_IO_110_mb1_FB1_BB0_IO_100,
    input wire        mb1_FA1_BA2_IO_111_mb1_FB1_BB0_IO_101,
    input wire        mb1_FA1_BA2_IO_112_mb1_FB1_BB0_IO_098,
    input wire        mb1_FA1_BA2_IO_113_mb1_FB1_BB0_IO_099,
    input wire        mb1_FA1_BA2_IO_114_mb1_FB1_BB0_IO_116,
    input wire        mb1_FA1_BA2_IO_115_mb1_FB1_BB0_IO_117,
    input wire        mb1_FA1_BA2_IO_116_mb1_FB1_BB0_IO_114,
    input wire        mb1_FA1_BA2_IO_117_mb1_FB1_BB0_IO_115,
    input wire        mb1_FA1_BA2_IO_118_mb1_FB1_BB0_IO_132,
    input wire        mb1_FA1_BA2_IO_119_mb1_FB1_BB0_IO_133,
    input wire        mb1_FA1_BA2_IO_120_mb1_FB1_BB0_IO_130,
    input wire        mb1_FA1_BA2_IO_121_mb1_FB1_BB0_IO_131,
    input wire        mb1_FA1_BA2_IO_122_mb1_FB1_BB0_IO_108,
    input wire        mb1_FA1_BA2_IO_123_mb1_FB1_BB0_IO_109,
    input wire        mb1_FA1_BA2_IO_124_mb1_FB1_BB0_IO_126,
    input wire        mb1_FA1_BA2_IO_125_mb1_FB1_BB0_IO_127,
    input wire        mb1_FA1_BA2_IO_126_mb1_FB1_BB0_IO_124,
    input wire        mb1_FA1_BA2_IO_127_mb1_FB1_BB0_IO_125,
    input wire        mb1_FA1_BA2_IO_130_mb1_FB1_BB0_IO_120,
    input wire        mb1_FA1_BA2_IO_131_mb1_FB1_BB0_IO_121,
    input wire        mb1_FA1_BA2_IO_132_mb1_FB1_BB0_IO_118,
    input wire        mb1_FA1_BA2_IO_133_mb1_FB1_BB0_IO_119,
    input wire        mb1_FA1_BA2_IO_134_mb1_FB1_BB0_IO_136,
    input wire        mb1_FA1_BA2_IO_136_mb1_FB1_BB0_IO_134,
    input wire        mb1_FA1_TB1_CLKIO_N_0_mb1_FB1_BB1_CLKIO_N_7,
    input wire        mb1_FA1_TB1_CLKIO_N_1_mb1_FB1_BB1_CLKIO_N_6,
    input wire        mb1_FA1_TB1_CLKIO_N_2_mb1_FB1_BB1_CLKIO_N_4,
    input wire        mb1_FA1_TB1_CLKIO_N_3_mb1_FB1_BB1_CLKIO_N_3,
    input wire        mb1_FA1_TB1_CLKIO_N_4_mb1_FB1_BB1_CLKIO_N_2,
    input wire        mb1_FA1_TB1_CLKIO_N_5_mb1_FB1_BB1_IO_010,
    input wire        mb1_FA1_TB1_CLKIO_N_6_mb1_FB1_BB1_CLKIO_N_1,
    input wire        mb1_FA1_TB1_CLKIO_N_7_mb1_FB1_BB1_CLKIO_N_0,
    input wire        mb1_FA1_TB1_CLKIO_P_0_mb1_FB1_BB1_CLKIO_P_7,
    input wire        mb1_FA1_TB1_CLKIO_P_1_mb1_FB1_BB1_CLKIO_P_6,
    input wire        mb1_FA1_TB1_CLKIO_P_2_mb1_FB1_BB1_CLKIO_P_4,
    input wire        mb1_FA1_TB1_CLKIO_P_3_mb1_FB1_BB1_CLKIO_P_3,
    input wire        mb1_FA1_TB1_CLKIO_P_4_mb1_FB1_BB1_CLKIO_P_2,
    input wire        mb1_FA1_TB1_CLKIO_P_5_mb1_FB1_BB1_IO_011,
    input wire        mb1_FA1_TB1_CLKIO_P_6_mb1_FB1_BB1_CLKIO_P_1,
    input wire        mb1_FA1_TB1_CLKIO_P_7_mb1_FB1_BB1_CLKIO_P_0,
    input wire        mb1_FA1_TB1_IO_004_mb1_FB1_BB1_IO_006,
    input wire        mb1_FA1_TB1_IO_005_mb1_FB1_BB1_IO_007,
    input wire        mb1_FA1_TB1_IO_006_mb1_FB1_BB1_IO_004,
    input wire        mb1_FA1_TB1_IO_007_mb1_FB1_BB1_IO_005,
    input wire        mb1_FA1_TB1_IO_008_mb1_FB1_BB1_IO_022,
    input wire        mb1_FA1_TB1_IO_009_mb1_FB1_BB1_IO_023,
    input wire        mb1_FA1_TB1_IO_010_mb1_FB1_BB1_CLKIO_N_5,
    input wire        mb1_FA1_TB1_IO_011_mb1_FB1_BB1_CLKIO_P_5,
    input wire        mb1_FA1_TB1_IO_012_mb1_FB1_BB1_IO_012,
    input wire        mb1_FA1_TB1_IO_013_mb1_FB1_BB1_IO_013,
    input wire        mb1_FA1_TB1_IO_014_mb1_FB1_BB1_IO_016,
    input wire        mb1_FA1_TB1_IO_015_mb1_FB1_BB1_IO_017,
    input wire        mb1_FA1_TB1_IO_016_mb1_FB1_BB1_IO_014,
    input wire        mb1_FA1_TB1_IO_017_mb1_FB1_BB1_IO_015,
    input wire        mb1_FA1_TB1_IO_018_mb1_FB1_BB1_IO_032,
    input wire        mb1_FA1_TB1_IO_019_mb1_FB1_BB1_IO_033,
    input wire        mb1_FA1_TB1_IO_020_mb1_FB1_BB1_IO_030,
    input wire        mb1_FA1_TB1_IO_021_mb1_FB1_BB1_IO_031,
    input wire        mb1_FA1_TB1_IO_022_mb1_FB1_BB1_IO_008,
    input wire        mb1_FA1_TB1_IO_023_mb1_FB1_BB1_IO_009,
    input wire        mb1_FA1_TB1_IO_024_mb1_FB1_BB1_IO_026,
    input wire        mb1_FA1_TB1_IO_025_mb1_FB1_BB1_IO_027,
    input wire        mb1_FA1_TB1_IO_026_mb1_FB1_BB1_IO_024,
    input wire        mb1_FA1_TB1_IO_027_mb1_FB1_BB1_IO_025,
    input wire        mb1_FA1_TB1_IO_028_mb1_FB1_BB1_IO_042,
    input wire        mb1_FA1_TB1_IO_029_mb1_FB1_BB1_IO_043,
    input wire        mb1_FA1_TB1_IO_030_mb1_FB1_BB1_IO_020,
    input wire        mb1_FA1_TB1_IO_031_mb1_FB1_BB1_IO_021,
    input wire        mb1_FA1_TB1_IO_032_mb1_FB1_BB1_IO_018,
    input wire        mb1_FA1_TB1_IO_033_mb1_FB1_BB1_IO_019,
    input wire        mb1_FA1_TB1_IO_034_mb1_FB1_BB1_IO_036,
    input wire        mb1_FA1_TB1_IO_035_mb1_FB1_BB1_IO_037,
    input wire        mb1_FA1_TB1_IO_036_mb1_FB1_BB1_IO_034,
    input wire        mb1_FA1_TB1_IO_037_mb1_FB1_BB1_IO_035,
    input wire        mb1_FA1_TB1_IO_038_mb1_FB1_BB1_IO_052,
    input wire        mb1_FA1_TB1_IO_039_mb1_FB1_BB1_IO_053,
    input wire        mb1_FA1_TB1_IO_040_mb1_FB1_BB1_IO_050,
    input wire        mb1_FA1_TB1_IO_041_mb1_FB1_BB1_IO_051,
    input wire        mb1_FA1_TB1_IO_042_mb1_FB1_BB1_IO_028,
    input wire        mb1_FA1_TB1_IO_043_mb1_FB1_BB1_IO_029,
    input wire        mb1_FA1_TB1_IO_044_mb1_FB1_BB1_IO_046,
    input wire        mb1_FA1_TB1_IO_045_mb1_FB1_BB1_IO_047,
    input wire        mb1_FA1_TB1_IO_046_mb1_FB1_BB1_IO_044,
    input wire        mb1_FA1_TB1_IO_047_mb1_FB1_BB1_IO_045,
    input wire        mb1_FA1_TB1_IO_048_mb1_FB1_BB1_IO_062,
    input wire        mb1_FA1_TB1_IO_049_mb1_FB1_BB1_IO_063,
    input wire        mb1_FA1_TB1_IO_050_mb1_FB1_BB1_IO_040,
    input wire        mb1_FA1_TB1_IO_051_mb1_FB1_BB1_IO_041,
    input wire        mb1_FA1_TB1_IO_052_mb1_FB1_BB1_IO_038,
    input wire        mb1_FA1_TB1_IO_053_mb1_FB1_BB1_IO_039,
    input wire        mb1_FA1_TB1_IO_054_mb1_FB1_BB1_IO_056,
    input wire        mb1_FA1_TB1_IO_055_mb1_FB1_BB1_IO_057,
    input wire        mb1_FA1_TB1_IO_056_mb1_FB1_BB1_IO_054,
    input wire        mb1_FA1_TB1_IO_057_mb1_FB1_BB1_IO_055,
    input wire        mb1_FA1_TB1_IO_058_mb1_FB1_BB1_IO_072,
    input wire        mb1_FA1_TB1_IO_059_mb1_FB1_BB1_IO_073,
    input wire        mb1_FA1_TB1_IO_060_mb1_FB1_BB1_IO_070,
    input wire        mb1_FA1_TB1_IO_061_mb1_FB1_BB1_IO_071,
    input wire        mb1_FA1_TB1_IO_062_mb1_FB1_BB1_IO_048,
    input wire        mb1_FA1_TB1_IO_063_mb1_FB1_BB1_IO_049,
    input wire        mb1_FA1_TB1_IO_064_mb1_FB1_BB1_IO_066,
    input wire        mb1_FA1_TB1_IO_065_mb1_FB1_BB1_IO_067,
    input wire        mb1_FA1_TB1_IO_066_mb1_FB1_BB1_IO_064,
    input wire        mb1_FA1_TB1_IO_067_mb1_FB1_BB1_IO_065,
    input wire        mb1_FA1_TB1_IO_068_mb1_FB1_BB1_IO_082,
    input wire        mb1_FA1_TB1_IO_069_mb1_FB1_BB1_IO_083,
    input wire        mb1_FA1_TB1_IO_070_mb1_FB1_BB1_IO_060,
    input wire        mb1_FA1_TB1_IO_071_mb1_FB1_BB1_IO_061,
    input wire        mb1_FA1_TB1_IO_072_mb1_FB1_BB1_IO_058,
    input wire        mb1_FA1_TB1_IO_073_mb1_FB1_BB1_IO_059,
    input wire        mb1_FA1_TB1_IO_074_mb1_FB1_BB1_IO_076,
    input wire        mb1_FA1_TB1_IO_075_mb1_FB1_BB1_IO_077,
    input wire        mb1_FA1_TB1_IO_076_mb1_FB1_BB1_IO_074,
    input wire        mb1_FA1_TB1_IO_077_mb1_FB1_BB1_IO_075,
    input wire        mb1_FA1_TB1_IO_078_mb1_FB1_BB1_IO_092,
    input wire        mb1_FA1_TB1_IO_079_mb1_FB1_BB1_IO_093,
    input wire        mb1_FA1_TB1_IO_080_mb1_FB1_BB1_IO_090,
    input wire        mb1_FA1_TB1_IO_081_mb1_FB1_BB1_IO_091,
    input wire        mb1_FA1_TB1_IO_082_mb1_FB1_BB1_IO_068,
    input wire        mb1_FA1_TB1_IO_083_mb1_FB1_BB1_IO_069,
    input wire        mb1_FA1_TB1_IO_084_mb1_FB1_BB1_IO_086,
    input wire        mb1_FA1_TB1_IO_085_mb1_FB1_BB1_IO_087,
    input wire        mb1_FA1_TB1_IO_086_mb1_FB1_BB1_IO_084,
    input wire        mb1_FA1_TB1_IO_087_mb1_FB1_BB1_IO_085,
    input wire        mb1_FA1_TB1_IO_088_mb1_FB1_BB1_IO_102,
    input wire        mb1_FA1_TB1_IO_089_mb1_FB1_BB1_IO_103,
    input wire        mb1_FA1_TB1_IO_090_mb1_FB1_BB1_IO_080,
    input wire        mb1_FA1_TB1_IO_091_mb1_FB1_BB1_IO_081,
    input wire        mb1_FA1_TB1_IO_092_mb1_FB1_BB1_IO_078,
    input wire        mb1_FA1_TB1_IO_093_mb1_FB1_BB1_IO_079,
    input wire        mb1_FA1_TB1_IO_094_mb1_FB1_BB1_IO_096,
    input wire        mb1_FA1_TB1_IO_095_mb1_FB1_BB1_IO_097,
    input wire        mb1_FA1_TB1_IO_096_mb1_FB1_BB1_IO_094,
    input wire        mb1_FA1_TB1_IO_097_mb1_FB1_BB1_IO_095,
    input wire        mb1_FA1_TB1_IO_098_mb1_FB1_BB1_IO_112,
    input wire        mb1_FA1_TB1_IO_099_mb1_FB1_BB1_IO_113,
    input wire        mb1_FA1_TB1_IO_100_mb1_FB1_BB1_IO_110,
    input wire        mb1_FA1_TB1_IO_101_mb1_FB1_BB1_IO_111,
    input wire        mb1_FA1_TB1_IO_102_mb1_FB1_BB1_IO_088,
    input wire        mb1_FA1_TB1_IO_103_mb1_FB1_BB1_IO_089,
    input wire        mb1_FA1_TB1_IO_104_mb1_FB1_BB1_IO_106,
    input wire        mb1_FA1_TB1_IO_105_mb1_FB1_BB1_IO_107,
    input wire        mb1_FA1_TB1_IO_106_mb1_FB1_BB1_IO_104,
    input wire        mb1_FA1_TB1_IO_107_mb1_FB1_BB1_IO_105,
    input wire        mb1_FA1_TB1_IO_108_mb1_FB1_BB1_IO_122,
    input wire        mb1_FA1_TB1_IO_109_mb1_FB1_BB1_IO_123,
    input wire        mb1_FA1_TB1_IO_110_mb1_FB1_BB1_IO_100,
    input wire        mb1_FA1_TB1_IO_111_mb1_FB1_BB1_IO_101,
    input wire        mb1_FA1_TB1_IO_112_mb1_FB1_BB1_IO_098,
    input wire        mb1_FA1_TB1_IO_113_mb1_FB1_BB1_IO_099,
    input wire        mb1_FA1_TB1_IO_114_mb1_FB1_BB1_IO_116,
    input wire        mb1_FA1_TB1_IO_115_mb1_FB1_BB1_IO_117,
    input wire        mb1_FA1_TB1_IO_116_mb1_FB1_BB1_IO_114,
    input wire        mb1_FA1_TB1_IO_117_mb1_FB1_BB1_IO_115,
    input wire        mb1_FA1_TB1_IO_118_mb1_FB1_BB1_IO_132,
    input wire        mb1_FA1_TB1_IO_119_mb1_FB1_BB1_IO_133,
    input wire        mb1_FA1_TB1_IO_120_mb1_FB1_BB1_IO_130,
    input wire        mb1_FA1_TB1_IO_121_mb1_FB1_BB1_IO_131,
    input wire        mb1_FA1_TB1_IO_122_mb1_FB1_BB1_IO_108,
    input wire        mb1_FA1_TB1_IO_123_mb1_FB1_BB1_IO_109,
    input wire        mb1_FA1_TB1_IO_124_mb1_FB1_BB1_IO_126,
    input wire        mb1_FA1_TB1_IO_125_mb1_FB1_BB1_IO_127,
    input wire        mb1_FA1_TB1_IO_126_mb1_FB1_BB1_IO_124,
    input wire        mb1_FA1_TB1_IO_127_mb1_FB1_BB1_IO_125,
    input wire        mb1_FA1_TB1_IO_130_mb1_FB1_BB1_IO_120,
    input wire        mb1_FA1_TB1_IO_131_mb1_FB1_BB1_IO_121,
    input wire        mb1_FA1_TB1_IO_132_mb1_FB1_BB1_IO_118,
    input wire        mb1_FA1_TB1_IO_133_mb1_FB1_BB1_IO_119,
    input wire        mb1_FA1_TB1_IO_134_mb1_FB1_BB1_IO_136,
    input wire        mb1_FA1_TB1_IO_136_mb1_FB1_BB1_IO_134,
    input wire        mb1_FA1_BB0_CLKIO_N_0_mb1_FB1_BB2_CLKIO_N_7,
    input wire        mb1_FA1_BB0_CLKIO_N_1_mb1_FB1_BB2_CLKIO_N_6,
    input wire        mb1_FA1_BB0_CLKIO_N_2_mb1_FB1_BB2_CLKIO_N_4,
    input wire        mb1_FA1_BB0_CLKIO_N_3_mb1_FB1_BB2_CLKIO_N_3,
    input wire        mb1_FA1_BB0_CLKIO_N_4_mb1_FB1_BB2_CLKIO_N_2,
    input wire        mb1_FA1_BB0_CLKIO_N_5_mb1_FB1_BB2_IO_010,
    input wire        mb1_FA1_BB0_CLKIO_N_6_mb1_FB1_BB2_CLKIO_N_1,
    input wire        mb1_FA1_BB0_CLKIO_N_7_mb1_FB1_BB2_CLKIO_N_0,
    input wire        mb1_FA1_BB0_CLKIO_P_0_mb1_FB1_BB2_CLKIO_P_7,
    input wire        mb1_FA1_BB0_CLKIO_P_1_mb1_FB1_BB2_CLKIO_P_6,
    input wire        mb1_FA1_BB0_CLKIO_P_2_mb1_FB1_BB2_CLKIO_P_4,
    input wire        mb1_FA1_BB0_CLKIO_P_3_mb1_FB1_BB2_CLKIO_P_3,
    input wire        mb1_FA1_BB0_CLKIO_P_4_mb1_FB1_BB2_CLKIO_P_2,
    input wire        mb1_FA1_BB0_CLKIO_P_5_mb1_FB1_BB2_IO_011,
    input wire        mb1_FA1_BB0_CLKIO_P_6_mb1_FB1_BB2_CLKIO_P_1,
    input wire        mb1_FA1_BB0_CLKIO_P_7_mb1_FB1_BB2_CLKIO_P_0,
    input wire        mb1_FA1_BB0_IO_004_mb1_FB1_BB2_IO_006,
    input wire        mb1_FA1_BB0_IO_005_mb1_FB1_BB2_IO_007,
    input wire        mb1_FA1_BB0_IO_006_mb1_FB1_BB2_IO_004,
    input wire        mb1_FA1_BB0_IO_007_mb1_FB1_BB2_IO_005,
    input wire        mb1_FA1_BB0_IO_008_mb1_FB1_BB2_IO_022,
    input wire        mb1_FA1_BB0_IO_009_mb1_FB1_BB2_IO_023,
    input wire        mb1_FA1_BB0_IO_010_mb1_FB1_BB2_CLKIO_N_5,
    input wire        mb1_FA1_BB0_IO_011_mb1_FB1_BB2_CLKIO_P_5,
    input wire        mb1_FA1_BB0_IO_012_mb1_FB1_BB2_IO_012,
    input wire        mb1_FA1_BB0_IO_013_mb1_FB1_BB2_IO_013,
    input wire        mb1_FA1_BB0_IO_014_mb1_FB1_BB2_IO_016,
    input wire        mb1_FA1_BB0_IO_015_mb1_FB1_BB2_IO_017,
    input wire        mb1_FA1_BB0_IO_016_mb1_FB1_BB2_IO_014,
    input wire        mb1_FA1_BB0_IO_017_mb1_FB1_BB2_IO_015,
    input wire        mb1_FA1_BB0_IO_018_mb1_FB1_BB2_IO_032,
    input wire        mb1_FA1_BB0_IO_019_mb1_FB1_BB2_IO_033,
    input wire        mb1_FA1_BB0_IO_020_mb1_FB1_BB2_IO_030,
    input wire        mb1_FA1_BB0_IO_021_mb1_FB1_BB2_IO_031,
    input wire        mb1_FA1_BB0_IO_022_mb1_FB1_BB2_IO_008,
    input wire        mb1_FA1_BB0_IO_023_mb1_FB1_BB2_IO_009,
    input wire        mb1_FA1_BB0_IO_024_mb1_FB1_BB2_IO_026,
    input wire        mb1_FA1_BB0_IO_025_mb1_FB1_BB2_IO_027,
    input wire        mb1_FA1_BB0_IO_026_mb1_FB1_BB2_IO_024,
    input wire        mb1_FA1_BB0_IO_027_mb1_FB1_BB2_IO_025,
    input wire        mb1_FA1_BB0_IO_028_mb1_FB1_BB2_IO_042,
    input wire        mb1_FA1_BB0_IO_029_mb1_FB1_BB2_IO_043,
    input wire        mb1_FA1_BB0_IO_030_mb1_FB1_BB2_IO_020,
    input wire        mb1_FA1_BB0_IO_031_mb1_FB1_BB2_IO_021,
    input wire        mb1_FA1_BB0_IO_032_mb1_FB1_BB2_IO_018,
    input wire        mb1_FA1_BB0_IO_033_mb1_FB1_BB2_IO_019,
    input wire        mb1_FA1_BB0_IO_034_mb1_FB1_BB2_IO_036,
    input wire        mb1_FA1_BB0_IO_035_mb1_FB1_BB2_IO_037,
    input wire        mb1_FA1_BB0_IO_036_mb1_FB1_BB2_IO_034,
    input wire        mb1_FA1_BB0_IO_037_mb1_FB1_BB2_IO_035,
    input wire        mb1_FA1_BB0_IO_038_mb1_FB1_BB2_IO_052,
    input wire        mb1_FA1_BB0_IO_039_mb1_FB1_BB2_IO_053,
    input wire        mb1_FA1_BB0_IO_040_mb1_FB1_BB2_IO_050,
    input wire        mb1_FA1_BB0_IO_041_mb1_FB1_BB2_IO_051,
    input wire        mb1_FA1_BB0_IO_042_mb1_FB1_BB2_IO_028,
    input wire        mb1_FA1_BB0_IO_043_mb1_FB1_BB2_IO_029,
    input wire        mb1_FA1_BB0_IO_044_mb1_FB1_BB2_IO_046,
    input wire        mb1_FA1_BB0_IO_045_mb1_FB1_BB2_IO_047,
    input wire        mb1_FA1_BB0_IO_046_mb1_FB1_BB2_IO_044,
    input wire        mb1_FA1_BB0_IO_047_mb1_FB1_BB2_IO_045,
    input wire        mb1_FA1_BB0_IO_048_mb1_FB1_BB2_IO_062,
    input wire        mb1_FA1_BB0_IO_049_mb1_FB1_BB2_IO_063,
    input wire        mb1_FA1_BB0_IO_050_mb1_FB1_BB2_IO_040,
    input wire        mb1_FA1_BB0_IO_051_mb1_FB1_BB2_IO_041,
    input wire        mb1_FA1_BB0_IO_052_mb1_FB1_BB2_IO_038,
    input wire        mb1_FA1_BB0_IO_053_mb1_FB1_BB2_IO_039,
    input wire        mb1_FA1_BB0_IO_054_mb1_FB1_BB2_IO_056,
    input wire        mb1_FA1_BB0_IO_055_mb1_FB1_BB2_IO_057,
    input wire        mb1_FA1_BB0_IO_056_mb1_FB1_BB2_IO_054,
    input wire        mb1_FA1_BB0_IO_057_mb1_FB1_BB2_IO_055,
    input wire        mb1_FA1_BB0_IO_058_mb1_FB1_BB2_IO_072,
    input wire        mb1_FA1_BB0_IO_059_mb1_FB1_BB2_IO_073,
    input wire        mb1_FA1_BB0_IO_060_mb1_FB1_BB2_IO_070,
    input wire        mb1_FA1_BB0_IO_061_mb1_FB1_BB2_IO_071,
    input wire        mb1_FA1_BB0_IO_062_mb1_FB1_BB2_IO_048,
    input wire        mb1_FA1_BB0_IO_063_mb1_FB1_BB2_IO_049,
    input wire        mb1_FA1_BB0_IO_064_mb1_FB1_BB2_IO_066,
    input wire        mb1_FA1_BB0_IO_065_mb1_FB1_BB2_IO_067,
    input wire        mb1_FA1_BB0_IO_066_mb1_FB1_BB2_IO_064,
    input wire        mb1_FA1_BB0_IO_067_mb1_FB1_BB2_IO_065,
    input wire        mb1_FA1_BB0_IO_068_mb1_FB1_BB2_IO_082,
    input wire        mb1_FA1_BB0_IO_069_mb1_FB1_BB2_IO_083,
    input wire        mb1_FA1_BB0_IO_070_mb1_FB1_BB2_IO_060,
    input wire        mb1_FA1_BB0_IO_071_mb1_FB1_BB2_IO_061,
    input wire        mb1_FA1_BB0_IO_072_mb1_FB1_BB2_IO_058,
    input wire        mb1_FA1_BB0_IO_073_mb1_FB1_BB2_IO_059,
    input wire        mb1_FA1_BB0_IO_074_mb1_FB1_BB2_IO_076,
    input wire        mb1_FA1_BB0_IO_075_mb1_FB1_BB2_IO_077,
    input wire        mb1_FA1_BB0_IO_076_mb1_FB1_BB2_IO_074,
    input wire        mb1_FA1_BB0_IO_077_mb1_FB1_BB2_IO_075,
    input wire        mb1_FA1_BB0_IO_078_mb1_FB1_BB2_IO_092,
    input wire        mb1_FA1_BB0_IO_079_mb1_FB1_BB2_IO_093,
    input wire        mb1_FA1_BB0_IO_080_mb1_FB1_BB2_IO_090,
    input wire        mb1_FA1_BB0_IO_081_mb1_FB1_BB2_IO_091,
    input wire        mb1_FA1_BB0_IO_082_mb1_FB1_BB2_IO_068,
    input wire        mb1_FA1_BB0_IO_083_mb1_FB1_BB2_IO_069,
    input wire        mb1_FA1_BB0_IO_084_mb1_FB1_BB2_IO_086,
    input wire        mb1_FA1_BB0_IO_085_mb1_FB1_BB2_IO_087,
    input wire        mb1_FA1_BB0_IO_086_mb1_FB1_BB2_IO_084,
    input wire        mb1_FA1_BB0_IO_087_mb1_FB1_BB2_IO_085,
    input wire        mb1_FA1_BB0_IO_088_mb1_FB1_BB2_IO_102,
    input wire        mb1_FA1_BB0_IO_089_mb1_FB1_BB2_IO_103,
    input wire        mb1_FA1_BB0_IO_090_mb1_FB1_BB2_IO_080,
    input wire        mb1_FA1_BB0_IO_091_mb1_FB1_BB2_IO_081,
    input wire        mb1_FA1_BB0_IO_092_mb1_FB1_BB2_IO_078,
    input wire        mb1_FA1_BB0_IO_093_mb1_FB1_BB2_IO_079,
    input wire        mb1_FA1_BB0_IO_094_mb1_FB1_BB2_IO_096,
    input wire        mb1_FA1_BB0_IO_095_mb1_FB1_BB2_IO_097,
    input wire        mb1_FA1_BB0_IO_096_mb1_FB1_BB2_IO_094,
    input wire        mb1_FA1_BB0_IO_097_mb1_FB1_BB2_IO_095,
    input wire        mb1_FA1_BB0_IO_098_mb1_FB1_BB2_IO_112,
    input wire        mb1_FA1_BB0_IO_099_mb1_FB1_BB2_IO_113,
    input wire        mb1_FA1_BB0_IO_100_mb1_FB1_BB2_IO_110,
    input wire        mb1_FA1_BB0_IO_101_mb1_FB1_BB2_IO_111,
    input wire        mb1_FA1_BB0_IO_102_mb1_FB1_BB2_IO_088,
    input wire        mb1_FA1_BB0_IO_103_mb1_FB1_BB2_IO_089,
    input wire        mb1_FA1_BB0_IO_104_mb1_FB1_BB2_IO_106,
    input wire        mb1_FA1_BB0_IO_105_mb1_FB1_BB2_IO_107,
    input wire        mb1_FA1_BB0_IO_106_mb1_FB1_BB2_IO_104,
    input wire        mb1_FA1_BB0_IO_107_mb1_FB1_BB2_IO_105,
    input wire        mb1_FA1_BB0_IO_108_mb1_FB1_BB2_IO_122,
    input wire        mb1_FA1_BB0_IO_109_mb1_FB1_BB2_IO_123,
    input wire        mb1_FA1_BB0_IO_110_mb1_FB1_BB2_IO_100,
    input wire        mb1_FA1_BB0_IO_111_mb1_FB1_BB2_IO_101,
    input wire        mb1_FA1_BB0_IO_112_mb1_FB1_BB2_IO_098,
    input wire        mb1_FA1_BB0_IO_113_mb1_FB1_BB2_IO_099,
    input wire        mb1_FA1_BB0_IO_114_mb1_FB1_BB2_IO_116,
    input wire        mb1_FA1_BB0_IO_115_mb1_FB1_BB2_IO_117,
    input wire        mb1_FA1_BB0_IO_116_mb1_FB1_BB2_IO_114,
    input wire        mb1_FA1_BB0_IO_117_mb1_FB1_BB2_IO_115,
    input wire        mb1_FA1_BB0_IO_118_mb1_FB1_BB2_IO_132,
    input wire        mb1_FA1_BB0_IO_119_mb1_FB1_BB2_IO_133,
    input wire        mb1_FA1_BB0_IO_120_mb1_FB1_BB2_IO_130,
    input wire        mb1_FA1_BB0_IO_121_mb1_FB1_BB2_IO_131,
    input wire        mb1_FA1_BB0_IO_122_mb1_FB1_BB2_IO_108,
    input wire        mb1_FA1_BB0_IO_123_mb1_FB1_BB2_IO_109,
    input wire        mb1_FA1_BB0_IO_124_mb1_FB1_BB2_IO_126,
    input wire        mb1_FA1_BB0_IO_125_mb1_FB1_BB2_IO_127,
    input wire        mb1_FA1_BB0_IO_126_mb1_FB1_BB2_IO_124,
    input wire        mb1_FA1_BB0_IO_127_mb1_FB1_BB2_IO_125,
    input wire        mb1_FA1_BB0_IO_130_mb1_FB1_BB2_IO_120,
    input wire        mb1_FA1_BB0_IO_131_mb1_FB1_BB2_IO_121,
    input wire        mb1_FA1_BB0_IO_132_mb1_FB1_BB2_IO_118,
    input wire        mb1_FA1_BB0_IO_133_mb1_FB1_BB2_IO_119,
    input wire        mb1_FA1_BB0_IO_134_mb1_FB1_BB2_IO_136,
    input wire        mb1_FA1_BB0_IO_136_mb1_FB1_BB2_IO_134);

  localparam TX_PINS            = 730;
  localparam RX_PINS            = 876;
  localparam USE_CLK_INPUT_BUFG = 0;

  wire [RX_PINS-1:0] rx_pin;
  wire [TX_PINS-1:0] tx_pin;

  assign mb1_FB1_TA1_CLKIO_N_0_mb1_FB2_BB0_CLKIO_N_7 = tx_pin[0];
  assign mb1_FB1_TA1_CLKIO_N_1_mb1_FB2_BB0_CLKIO_N_6 = tx_pin[1];
  assign mb1_FB1_TA1_CLKIO_N_2_mb1_FB2_BB0_CLKIO_N_4 = tx_pin[2];
  assign mb1_FB1_TA1_CLKIO_N_3_mb1_FB2_BB0_CLKIO_N_3 = tx_pin[3];
  assign mb1_FB1_TA1_CLKIO_N_4_mb1_FB2_BB0_CLKIO_N_2 = tx_pin[4];
  assign mb1_FB1_TA1_CLKIO_N_5_mb1_FB2_BB0_IO_010 = tx_pin[5];
  assign mb1_FB1_TA1_CLKIO_N_6_mb1_FB2_BB0_CLKIO_N_1 = tx_pin[6];
  assign mb1_FB1_TA1_CLKIO_N_7_mb1_FB2_BB0_CLKIO_N_0 = tx_pin[7];
  assign mb1_FB1_TA1_CLKIO_P_0_mb1_FB2_BB0_CLKIO_P_7 = tx_pin[8];
  assign mb1_FB1_TA1_CLKIO_P_1_mb1_FB2_BB0_CLKIO_P_6 = tx_pin[9];
  assign mb1_FB1_TA1_CLKIO_P_2_mb1_FB2_BB0_CLKIO_P_4 = tx_pin[10];
  assign mb1_FB1_TA1_CLKIO_P_3_mb1_FB2_BB0_CLKIO_P_3 = tx_pin[11];
  assign mb1_FB1_TA1_CLKIO_P_4_mb1_FB2_BB0_CLKIO_P_2 = tx_pin[12];
  assign mb1_FB1_TA1_CLKIO_P_5_mb1_FB2_BB0_IO_011 = tx_pin[13];
  assign mb1_FB1_TA1_CLKIO_P_6_mb1_FB2_BB0_CLKIO_P_1 = tx_pin[14];
  assign mb1_FB1_TA1_CLKIO_P_7_mb1_FB2_BB0_CLKIO_P_0 = tx_pin[15];
  assign mb1_FB1_TA1_IO_004_mb1_FB2_BB0_IO_006 = tx_pin[16];
  assign mb1_FB1_TA1_IO_005_mb1_FB2_BB0_IO_007 = tx_pin[17];
  assign mb1_FB1_TA1_IO_006_mb1_FB2_BB0_IO_004 = tx_pin[18];
  assign mb1_FB1_TA1_IO_007_mb1_FB2_BB0_IO_005 = tx_pin[19];
  assign mb1_FB1_TA1_IO_008_mb1_FB2_BB0_IO_022 = tx_pin[20];
  assign mb1_FB1_TA1_IO_009_mb1_FB2_BB0_IO_023 = tx_pin[21];
  assign mb1_FB1_TA1_IO_010_mb1_FB2_BB0_CLKIO_N_5 = tx_pin[22];
  assign mb1_FB1_TA1_IO_011_mb1_FB2_BB0_CLKIO_P_5 = tx_pin[23];
  assign mb1_FB1_TA1_IO_012_mb1_FB2_BB0_IO_012 = tx_pin[24];
  assign mb1_FB1_TA1_IO_013_mb1_FB2_BB0_IO_013 = tx_pin[25];
  assign mb1_FB1_TA1_IO_014_mb1_FB2_BB0_IO_016 = tx_pin[26];
  assign mb1_FB1_TA1_IO_015_mb1_FB2_BB0_IO_017 = tx_pin[27];
  assign mb1_FB1_TA1_IO_016_mb1_FB2_BB0_IO_014 = tx_pin[28];
  assign mb1_FB1_TA1_IO_017_mb1_FB2_BB0_IO_015 = tx_pin[29];
  assign mb1_FB1_TA1_IO_018_mb1_FB2_BB0_IO_032 = tx_pin[30];
  assign mb1_FB1_TA1_IO_019_mb1_FB2_BB0_IO_033 = tx_pin[31];
  assign mb1_FB1_TA1_IO_020_mb1_FB2_BB0_IO_030 = tx_pin[32];
  assign mb1_FB1_TA1_IO_021_mb1_FB2_BB0_IO_031 = tx_pin[33];
  assign mb1_FB1_TA1_IO_022_mb1_FB2_BB0_IO_008 = tx_pin[34];
  assign mb1_FB1_TA1_IO_023_mb1_FB2_BB0_IO_009 = tx_pin[35];
  assign mb1_FB1_TA1_IO_024_mb1_FB2_BB0_IO_026 = tx_pin[36];
  assign mb1_FB1_TA1_IO_025_mb1_FB2_BB0_IO_027 = tx_pin[37];
  assign mb1_FB1_TA1_IO_026_mb1_FB2_BB0_IO_024 = tx_pin[38];
  assign mb1_FB1_TA1_IO_027_mb1_FB2_BB0_IO_025 = tx_pin[39];
  assign mb1_FB1_TA1_IO_028_mb1_FB2_BB0_IO_042 = tx_pin[40];
  assign mb1_FB1_TA1_IO_029_mb1_FB2_BB0_IO_043 = tx_pin[41];
  assign mb1_FB1_TA1_IO_030_mb1_FB2_BB0_IO_020 = tx_pin[42];
  assign mb1_FB1_TA1_IO_031_mb1_FB2_BB0_IO_021 = tx_pin[43];
  assign mb1_FB1_TA1_IO_032_mb1_FB2_BB0_IO_018 = tx_pin[44];
  assign mb1_FB1_TA1_IO_033_mb1_FB2_BB0_IO_019 = tx_pin[45];
  assign mb1_FB1_TA1_IO_034_mb1_FB2_BB0_IO_036 = tx_pin[46];
  assign mb1_FB1_TA1_IO_035_mb1_FB2_BB0_IO_037 = tx_pin[47];
  assign mb1_FB1_TA1_IO_036_mb1_FB2_BB0_IO_034 = tx_pin[48];
  assign mb1_FB1_TA1_IO_037_mb1_FB2_BB0_IO_035 = tx_pin[49];
  assign mb1_FB1_TA1_IO_038_mb1_FB2_BB0_IO_052 = tx_pin[50];
  assign mb1_FB1_TA1_IO_039_mb1_FB2_BB0_IO_053 = tx_pin[51];
  assign mb1_FB1_TA1_IO_040_mb1_FB2_BB0_IO_050 = tx_pin[52];
  assign mb1_FB1_TA1_IO_041_mb1_FB2_BB0_IO_051 = tx_pin[53];
  assign mb1_FB1_TA1_IO_042_mb1_FB2_BB0_IO_028 = tx_pin[54];
  assign mb1_FB1_TA1_IO_043_mb1_FB2_BB0_IO_029 = tx_pin[55];
  assign mb1_FB1_TA1_IO_044_mb1_FB2_BB0_IO_046 = tx_pin[56];
  assign mb1_FB1_TA1_IO_045_mb1_FB2_BB0_IO_047 = tx_pin[57];
  assign mb1_FB1_TA1_IO_046_mb1_FB2_BB0_IO_044 = tx_pin[58];
  assign mb1_FB1_TA1_IO_047_mb1_FB2_BB0_IO_045 = tx_pin[59];
  assign mb1_FB1_TA1_IO_048_mb1_FB2_BB0_IO_062 = tx_pin[60];
  assign mb1_FB1_TA1_IO_049_mb1_FB2_BB0_IO_063 = tx_pin[61];
  assign mb1_FB1_TA1_IO_050_mb1_FB2_BB0_IO_040 = tx_pin[62];
  assign mb1_FB1_TA1_IO_051_mb1_FB2_BB0_IO_041 = tx_pin[63];
  assign mb1_FB1_TA1_IO_052_mb1_FB2_BB0_IO_038 = tx_pin[64];
  assign mb1_FB1_TA1_IO_053_mb1_FB2_BB0_IO_039 = tx_pin[65];
  assign mb1_FB1_TA1_IO_054_mb1_FB2_BB0_IO_056 = tx_pin[66];
  assign mb1_FB1_TA1_IO_055_mb1_FB2_BB0_IO_057 = tx_pin[67];
  assign mb1_FB1_TA1_IO_056_mb1_FB2_BB0_IO_054 = tx_pin[68];
  assign mb1_FB1_TA1_IO_057_mb1_FB2_BB0_IO_055 = tx_pin[69];
  assign mb1_FB1_TA1_IO_058_mb1_FB2_BB0_IO_072 = tx_pin[70];
  assign mb1_FB1_TA1_IO_059_mb1_FB2_BB0_IO_073 = tx_pin[71];
  assign mb1_FB1_TA1_IO_060_mb1_FB2_BB0_IO_070 = tx_pin[72];
  assign mb1_FB1_TA1_IO_061_mb1_FB2_BB0_IO_071 = tx_pin[73];
  assign mb1_FB1_TA1_IO_062_mb1_FB2_BB0_IO_048 = tx_pin[74];
  assign mb1_FB1_TA1_IO_063_mb1_FB2_BB0_IO_049 = tx_pin[75];
  assign mb1_FB1_TA1_IO_064_mb1_FB2_BB0_IO_066 = tx_pin[76];
  assign mb1_FB1_TA1_IO_065_mb1_FB2_BB0_IO_067 = tx_pin[77];
  assign mb1_FB1_TA1_IO_066_mb1_FB2_BB0_IO_064 = tx_pin[78];
  assign mb1_FB1_TA1_IO_067_mb1_FB2_BB0_IO_065 = tx_pin[79];
  assign mb1_FB1_TA1_IO_068_mb1_FB2_BB0_IO_082 = tx_pin[80];
  assign mb1_FB1_TA1_IO_069_mb1_FB2_BB0_IO_083 = tx_pin[81];
  assign mb1_FB1_TA1_IO_070_mb1_FB2_BB0_IO_060 = tx_pin[82];
  assign mb1_FB1_TA1_IO_071_mb1_FB2_BB0_IO_061 = tx_pin[83];
  assign mb1_FB1_TA1_IO_072_mb1_FB2_BB0_IO_058 = tx_pin[84];
  assign mb1_FB1_TA1_IO_073_mb1_FB2_BB0_IO_059 = tx_pin[85];
  assign mb1_FB1_TA1_IO_074_mb1_FB2_BB0_IO_076 = tx_pin[86];
  assign mb1_FB1_TA1_IO_075_mb1_FB2_BB0_IO_077 = tx_pin[87];
  assign mb1_FB1_TA1_IO_076_mb1_FB2_BB0_IO_074 = tx_pin[88];
  assign mb1_FB1_TA1_IO_077_mb1_FB2_BB0_IO_075 = tx_pin[89];
  assign mb1_FB1_TA1_IO_078_mb1_FB2_BB0_IO_092 = tx_pin[90];
  assign mb1_FB1_TA1_IO_079_mb1_FB2_BB0_IO_093 = tx_pin[91];
  assign mb1_FB1_TA1_IO_080_mb1_FB2_BB0_IO_090 = tx_pin[92];
  assign mb1_FB1_TA1_IO_081_mb1_FB2_BB0_IO_091 = tx_pin[93];
  assign mb1_FB1_TA1_IO_082_mb1_FB2_BB0_IO_068 = tx_pin[94];
  assign mb1_FB1_TA1_IO_083_mb1_FB2_BB0_IO_069 = tx_pin[95];
  assign mb1_FB1_TA1_IO_084_mb1_FB2_BB0_IO_086 = tx_pin[96];
  assign mb1_FB1_TA1_IO_085_mb1_FB2_BB0_IO_087 = tx_pin[97];
  assign mb1_FB1_TA1_IO_086_mb1_FB2_BB0_IO_084 = tx_pin[98];
  assign mb1_FB1_TA1_IO_087_mb1_FB2_BB0_IO_085 = tx_pin[99];
  assign mb1_FB1_TA1_IO_088_mb1_FB2_BB0_IO_102 = tx_pin[100];
  assign mb1_FB1_TA1_IO_089_mb1_FB2_BB0_IO_103 = tx_pin[101];
  assign mb1_FB1_TA1_IO_090_mb1_FB2_BB0_IO_080 = tx_pin[102];
  assign mb1_FB1_TA1_IO_091_mb1_FB2_BB0_IO_081 = tx_pin[103];
  assign mb1_FB1_TA1_IO_092_mb1_FB2_BB0_IO_078 = tx_pin[104];
  assign mb1_FB1_TA1_IO_093_mb1_FB2_BB0_IO_079 = tx_pin[105];
  assign mb1_FB1_TA1_IO_094_mb1_FB2_BB0_IO_096 = tx_pin[106];
  assign mb1_FB1_TA1_IO_095_mb1_FB2_BB0_IO_097 = tx_pin[107];
  assign mb1_FB1_TA1_IO_096_mb1_FB2_BB0_IO_094 = tx_pin[108];
  assign mb1_FB1_TA1_IO_097_mb1_FB2_BB0_IO_095 = tx_pin[109];
  assign mb1_FB1_TA1_IO_098_mb1_FB2_BB0_IO_112 = tx_pin[110];
  assign mb1_FB1_TA1_IO_099_mb1_FB2_BB0_IO_113 = tx_pin[111];
  assign mb1_FB1_TA1_IO_100_mb1_FB2_BB0_IO_110 = tx_pin[112];
  assign mb1_FB1_TA1_IO_101_mb1_FB2_BB0_IO_111 = tx_pin[113];
  assign mb1_FB1_TA1_IO_102_mb1_FB2_BB0_IO_088 = tx_pin[114];
  assign mb1_FB1_TA1_IO_103_mb1_FB2_BB0_IO_089 = tx_pin[115];
  assign mb1_FB1_TA1_IO_104_mb1_FB2_BB0_IO_106 = tx_pin[116];
  assign mb1_FB1_TA1_IO_105_mb1_FB2_BB0_IO_107 = tx_pin[117];
  assign mb1_FB1_TA1_IO_106_mb1_FB2_BB0_IO_104 = tx_pin[118];
  assign mb1_FB1_TA1_IO_107_mb1_FB2_BB0_IO_105 = tx_pin[119];
  assign mb1_FB1_TA1_IO_108_mb1_FB2_BB0_IO_122 = tx_pin[120];
  assign mb1_FB1_TA1_IO_109_mb1_FB2_BB0_IO_123 = tx_pin[121];
  assign mb1_FB1_TA1_IO_110_mb1_FB2_BB0_IO_100 = tx_pin[122];
  assign mb1_FB1_TA1_IO_111_mb1_FB2_BB0_IO_101 = tx_pin[123];
  assign mb1_FB1_TA1_IO_112_mb1_FB2_BB0_IO_098 = tx_pin[124];
  assign mb1_FB1_TA1_IO_113_mb1_FB2_BB0_IO_099 = tx_pin[125];
  assign mb1_FB1_TA1_IO_114_mb1_FB2_BB0_IO_116 = tx_pin[126];
  assign mb1_FB1_TA1_IO_115_mb1_FB2_BB0_IO_117 = tx_pin[127];
  assign mb1_FB1_TA1_IO_116_mb1_FB2_BB0_IO_114 = tx_pin[128];
  assign mb1_FB1_TA1_IO_117_mb1_FB2_BB0_IO_115 = tx_pin[129];
  assign mb1_FB1_TA1_IO_118_mb1_FB2_BB0_IO_132 = tx_pin[130];
  assign mb1_FB1_TA1_IO_119_mb1_FB2_BB0_IO_133 = tx_pin[131];
  assign mb1_FB1_TA1_IO_120_mb1_FB2_BB0_IO_130 = tx_pin[132];
  assign mb1_FB1_TA1_IO_121_mb1_FB2_BB0_IO_131 = tx_pin[133];
  assign mb1_FB1_TA1_IO_122_mb1_FB2_BB0_IO_108 = tx_pin[134];
  assign mb1_FB1_TA1_IO_123_mb1_FB2_BB0_IO_109 = tx_pin[135];
  assign mb1_FB1_TA1_IO_124_mb1_FB2_BB0_IO_126 = tx_pin[136];
  assign mb1_FB1_TA1_IO_125_mb1_FB2_BB0_IO_127 = tx_pin[137];
  assign mb1_FB1_TA1_IO_126_mb1_FB2_BB0_IO_124 = tx_pin[138];
  assign mb1_FB1_TA1_IO_127_mb1_FB2_BB0_IO_125 = tx_pin[139];
  assign mb1_FB1_TA1_IO_130_mb1_FB2_BB0_IO_120 = tx_pin[140];
  assign mb1_FB1_TA1_IO_131_mb1_FB2_BB0_IO_121 = tx_pin[141];
  assign mb1_FB1_TA1_IO_132_mb1_FB2_BB0_IO_118 = tx_pin[142];
  assign mb1_FB1_TA1_IO_133_mb1_FB2_BB0_IO_119 = tx_pin[143];
  assign mb1_FB1_TA1_IO_134_mb1_FB2_BB0_IO_136 = tx_pin[144];
  assign mb1_FB1_TA1_IO_136_mb1_FB2_BB0_IO_134 = tx_pin[145];
  assign rx_pin[0] = mb1_FA1_TA1_CLKIO_N_0_mb1_FB1_TA2_CLKIO_N_7;
  assign rx_pin[1] = mb1_FA1_TA1_CLKIO_N_1_mb1_FB1_TA2_CLKIO_N_6;
  assign rx_pin[2] = mb1_FA1_TA1_CLKIO_N_2_mb1_FB1_TA2_CLKIO_N_4;
  assign rx_pin[3] = mb1_FA1_TA1_CLKIO_N_3_mb1_FB1_TA2_CLKIO_N_3;
  assign rx_pin[4] = mb1_FA1_TA1_CLKIO_N_4_mb1_FB1_TA2_CLKIO_N_2;
  assign rx_pin[5] = mb1_FA1_TA1_CLKIO_N_5_mb1_FB1_TA2_IO_010;
  assign rx_pin[6] = mb1_FA1_TA1_CLKIO_N_6_mb1_FB1_TA2_CLKIO_N_1;
  assign rx_pin[7] = mb1_FA1_TA1_CLKIO_N_7_mb1_FB1_TA2_CLKIO_N_0;
  assign rx_pin[8] = mb1_FA1_TA1_CLKIO_P_0_mb1_FB1_TA2_CLKIO_P_7;
  assign rx_pin[9] = mb1_FA1_TA1_CLKIO_P_1_mb1_FB1_TA2_CLKIO_P_6;
  assign rx_pin[10] = mb1_FA1_TA1_CLKIO_P_2_mb1_FB1_TA2_CLKIO_P_4;
  assign rx_pin[11] = mb1_FA1_TA1_CLKIO_P_3_mb1_FB1_TA2_CLKIO_P_3;
  assign rx_pin[12] = mb1_FA1_TA1_CLKIO_P_4_mb1_FB1_TA2_CLKIO_P_2;
  assign rx_pin[13] = mb1_FA1_TA1_CLKIO_P_5_mb1_FB1_TA2_IO_011;
  assign rx_pin[14] = mb1_FA1_TA1_CLKIO_P_6_mb1_FB1_TA2_CLKIO_P_1;
  assign rx_pin[15] = mb1_FA1_TA1_CLKIO_P_7_mb1_FB1_TA2_CLKIO_P_0;
  assign rx_pin[16] = mb1_FA1_TA1_IO_004_mb1_FB1_TA2_IO_006;
  assign rx_pin[17] = mb1_FA1_TA1_IO_005_mb1_FB1_TA2_IO_007;
  assign rx_pin[18] = mb1_FA1_TA1_IO_006_mb1_FB1_TA2_IO_004;
  assign rx_pin[19] = mb1_FA1_TA1_IO_007_mb1_FB1_TA2_IO_005;
  assign rx_pin[20] = mb1_FA1_TA1_IO_008_mb1_FB1_TA2_IO_022;
  assign rx_pin[21] = mb1_FA1_TA1_IO_009_mb1_FB1_TA2_IO_023;
  assign rx_pin[22] = mb1_FA1_TA1_IO_010_mb1_FB1_TA2_CLKIO_N_5;
  assign rx_pin[23] = mb1_FA1_TA1_IO_011_mb1_FB1_TA2_CLKIO_P_5;
  assign rx_pin[24] = mb1_FA1_TA1_IO_012_mb1_FB1_TA2_IO_012;
  assign rx_pin[25] = mb1_FA1_TA1_IO_013_mb1_FB1_TA2_IO_013;
  assign rx_pin[26] = mb1_FA1_TA1_IO_014_mb1_FB1_TA2_IO_016;
  assign rx_pin[27] = mb1_FA1_TA1_IO_015_mb1_FB1_TA2_IO_017;
  assign rx_pin[28] = mb1_FA1_TA1_IO_016_mb1_FB1_TA2_IO_014;
  assign rx_pin[29] = mb1_FA1_TA1_IO_017_mb1_FB1_TA2_IO_015;
  assign rx_pin[30] = mb1_FA1_TA1_IO_018_mb1_FB1_TA2_IO_032;
  assign rx_pin[31] = mb1_FA1_TA1_IO_019_mb1_FB1_TA2_IO_033;
  assign rx_pin[32] = mb1_FA1_TA1_IO_020_mb1_FB1_TA2_IO_030;
  assign rx_pin[33] = mb1_FA1_TA1_IO_021_mb1_FB1_TA2_IO_031;
  assign rx_pin[34] = mb1_FA1_TA1_IO_022_mb1_FB1_TA2_IO_008;
  assign rx_pin[35] = mb1_FA1_TA1_IO_023_mb1_FB1_TA2_IO_009;
  assign rx_pin[36] = mb1_FA1_TA1_IO_024_mb1_FB1_TA2_IO_026;
  assign rx_pin[37] = mb1_FA1_TA1_IO_025_mb1_FB1_TA2_IO_027;
  assign rx_pin[38] = mb1_FA1_TA1_IO_026_mb1_FB1_TA2_IO_024;
  assign rx_pin[39] = mb1_FA1_TA1_IO_027_mb1_FB1_TA2_IO_025;
  assign rx_pin[40] = mb1_FA1_TA1_IO_028_mb1_FB1_TA2_IO_042;
  assign rx_pin[41] = mb1_FA1_TA1_IO_029_mb1_FB1_TA2_IO_043;
  assign rx_pin[42] = mb1_FA1_TA1_IO_030_mb1_FB1_TA2_IO_020;
  assign rx_pin[43] = mb1_FA1_TA1_IO_031_mb1_FB1_TA2_IO_021;
  assign rx_pin[44] = mb1_FA1_TA1_IO_032_mb1_FB1_TA2_IO_018;
  assign rx_pin[45] = mb1_FA1_TA1_IO_033_mb1_FB1_TA2_IO_019;
  assign rx_pin[46] = mb1_FA1_TA1_IO_034_mb1_FB1_TA2_IO_036;
  assign rx_pin[47] = mb1_FA1_TA1_IO_035_mb1_FB1_TA2_IO_037;
  assign rx_pin[48] = mb1_FA1_TA1_IO_036_mb1_FB1_TA2_IO_034;
  assign rx_pin[49] = mb1_FA1_TA1_IO_037_mb1_FB1_TA2_IO_035;
  assign rx_pin[50] = mb1_FA1_TA1_IO_038_mb1_FB1_TA2_IO_052;
  assign rx_pin[51] = mb1_FA1_TA1_IO_039_mb1_FB1_TA2_IO_053;
  assign rx_pin[52] = mb1_FA1_TA1_IO_040_mb1_FB1_TA2_IO_050;
  assign rx_pin[53] = mb1_FA1_TA1_IO_041_mb1_FB1_TA2_IO_051;
  assign rx_pin[54] = mb1_FA1_TA1_IO_042_mb1_FB1_TA2_IO_028;
  assign rx_pin[55] = mb1_FA1_TA1_IO_043_mb1_FB1_TA2_IO_029;
  assign rx_pin[56] = mb1_FA1_TA1_IO_044_mb1_FB1_TA2_IO_046;
  assign rx_pin[57] = mb1_FA1_TA1_IO_045_mb1_FB1_TA2_IO_047;
  assign rx_pin[58] = mb1_FA1_TA1_IO_046_mb1_FB1_TA2_IO_044;
  assign rx_pin[59] = mb1_FA1_TA1_IO_047_mb1_FB1_TA2_IO_045;
  assign rx_pin[60] = mb1_FA1_TA1_IO_048_mb1_FB1_TA2_IO_062;
  assign rx_pin[61] = mb1_FA1_TA1_IO_049_mb1_FB1_TA2_IO_063;
  assign rx_pin[62] = mb1_FA1_TA1_IO_050_mb1_FB1_TA2_IO_040;
  assign rx_pin[63] = mb1_FA1_TA1_IO_051_mb1_FB1_TA2_IO_041;
  assign rx_pin[64] = mb1_FA1_TA1_IO_052_mb1_FB1_TA2_IO_038;
  assign rx_pin[65] = mb1_FA1_TA1_IO_053_mb1_FB1_TA2_IO_039;
  assign rx_pin[66] = mb1_FA1_TA1_IO_054_mb1_FB1_TA2_IO_056;
  assign rx_pin[67] = mb1_FA1_TA1_IO_055_mb1_FB1_TA2_IO_057;
  assign rx_pin[68] = mb1_FA1_TA1_IO_056_mb1_FB1_TA2_IO_054;
  assign rx_pin[69] = mb1_FA1_TA1_IO_057_mb1_FB1_TA2_IO_055;
  assign rx_pin[70] = mb1_FA1_TA1_IO_058_mb1_FB1_TA2_IO_072;
  assign rx_pin[71] = mb1_FA1_TA1_IO_059_mb1_FB1_TA2_IO_073;
  assign rx_pin[72] = mb1_FA1_TA1_IO_060_mb1_FB1_TA2_IO_070;
  assign rx_pin[73] = mb1_FA1_TA1_IO_061_mb1_FB1_TA2_IO_071;
  assign rx_pin[74] = mb1_FA1_TA1_IO_062_mb1_FB1_TA2_IO_048;
  assign rx_pin[75] = mb1_FA1_TA1_IO_063_mb1_FB1_TA2_IO_049;
  assign rx_pin[76] = mb1_FA1_TA1_IO_064_mb1_FB1_TA2_IO_066;
  assign rx_pin[77] = mb1_FA1_TA1_IO_065_mb1_FB1_TA2_IO_067;
  assign rx_pin[78] = mb1_FA1_TA1_IO_066_mb1_FB1_TA2_IO_064;
  assign rx_pin[79] = mb1_FA1_TA1_IO_067_mb1_FB1_TA2_IO_065;
  assign rx_pin[80] = mb1_FA1_TA1_IO_068_mb1_FB1_TA2_IO_082;
  assign rx_pin[81] = mb1_FA1_TA1_IO_069_mb1_FB1_TA2_IO_083;
  assign rx_pin[82] = mb1_FA1_TA1_IO_070_mb1_FB1_TA2_IO_060;
  assign rx_pin[83] = mb1_FA1_TA1_IO_071_mb1_FB1_TA2_IO_061;
  assign rx_pin[84] = mb1_FA1_TA1_IO_072_mb1_FB1_TA2_IO_058;
  assign rx_pin[85] = mb1_FA1_TA1_IO_073_mb1_FB1_TA2_IO_059;
  assign rx_pin[86] = mb1_FA1_TA1_IO_074_mb1_FB1_TA2_IO_076;
  assign rx_pin[87] = mb1_FA1_TA1_IO_075_mb1_FB1_TA2_IO_077;
  assign rx_pin[88] = mb1_FA1_TA1_IO_076_mb1_FB1_TA2_IO_074;
  assign rx_pin[89] = mb1_FA1_TA1_IO_077_mb1_FB1_TA2_IO_075;
  assign rx_pin[90] = mb1_FA1_TA1_IO_078_mb1_FB1_TA2_IO_092;
  assign rx_pin[91] = mb1_FA1_TA1_IO_079_mb1_FB1_TA2_IO_093;
  assign rx_pin[92] = mb1_FA1_TA1_IO_080_mb1_FB1_TA2_IO_090;
  assign rx_pin[93] = mb1_FA1_TA1_IO_081_mb1_FB1_TA2_IO_091;
  assign rx_pin[94] = mb1_FA1_TA1_IO_082_mb1_FB1_TA2_IO_068;
  assign rx_pin[95] = mb1_FA1_TA1_IO_083_mb1_FB1_TA2_IO_069;
  assign rx_pin[96] = mb1_FA1_TA1_IO_084_mb1_FB1_TA2_IO_086;
  assign rx_pin[97] = mb1_FA1_TA1_IO_085_mb1_FB1_TA2_IO_087;
  assign rx_pin[98] = mb1_FA1_TA1_IO_086_mb1_FB1_TA2_IO_084;
  assign rx_pin[99] = mb1_FA1_TA1_IO_087_mb1_FB1_TA2_IO_085;
  assign rx_pin[100] = mb1_FA1_TA1_IO_088_mb1_FB1_TA2_IO_102;
  assign rx_pin[101] = mb1_FA1_TA1_IO_089_mb1_FB1_TA2_IO_103;
  assign rx_pin[102] = mb1_FA1_TA1_IO_090_mb1_FB1_TA2_IO_080;
  assign rx_pin[103] = mb1_FA1_TA1_IO_091_mb1_FB1_TA2_IO_081;
  assign rx_pin[104] = mb1_FA1_TA1_IO_092_mb1_FB1_TA2_IO_078;
  assign rx_pin[105] = mb1_FA1_TA1_IO_093_mb1_FB1_TA2_IO_079;
  assign rx_pin[106] = mb1_FA1_TA1_IO_094_mb1_FB1_TA2_IO_096;
  assign rx_pin[107] = mb1_FA1_TA1_IO_095_mb1_FB1_TA2_IO_097;
  assign rx_pin[108] = mb1_FA1_TA1_IO_096_mb1_FB1_TA2_IO_094;
  assign rx_pin[109] = mb1_FA1_TA1_IO_097_mb1_FB1_TA2_IO_095;
  assign rx_pin[110] = mb1_FA1_TA1_IO_098_mb1_FB1_TA2_IO_112;
  assign rx_pin[111] = mb1_FA1_TA1_IO_099_mb1_FB1_TA2_IO_113;
  assign rx_pin[112] = mb1_FA1_TA1_IO_100_mb1_FB1_TA2_IO_110;
  assign rx_pin[113] = mb1_FA1_TA1_IO_101_mb1_FB1_TA2_IO_111;
  assign rx_pin[114] = mb1_FA1_TA1_IO_102_mb1_FB1_TA2_IO_088;
  assign rx_pin[115] = mb1_FA1_TA1_IO_103_mb1_FB1_TA2_IO_089;
  assign rx_pin[116] = mb1_FA1_TA1_IO_104_mb1_FB1_TA2_IO_106;
  assign rx_pin[117] = mb1_FA1_TA1_IO_105_mb1_FB1_TA2_IO_107;
  assign rx_pin[118] = mb1_FA1_TA1_IO_106_mb1_FB1_TA2_IO_104;
  assign rx_pin[119] = mb1_FA1_TA1_IO_107_mb1_FB1_TA2_IO_105;
  assign rx_pin[120] = mb1_FA1_TA1_IO_108_mb1_FB1_TA2_IO_122;
  assign rx_pin[121] = mb1_FA1_TA1_IO_109_mb1_FB1_TA2_IO_123;
  assign rx_pin[122] = mb1_FA1_TA1_IO_110_mb1_FB1_TA2_IO_100;
  assign rx_pin[123] = mb1_FA1_TA1_IO_111_mb1_FB1_TA2_IO_101;
  assign rx_pin[124] = mb1_FA1_TA1_IO_112_mb1_FB1_TA2_IO_098;
  assign rx_pin[125] = mb1_FA1_TA1_IO_113_mb1_FB1_TA2_IO_099;
  assign rx_pin[126] = mb1_FA1_TA1_IO_114_mb1_FB1_TA2_IO_116;
  assign rx_pin[127] = mb1_FA1_TA1_IO_115_mb1_FB1_TA2_IO_117;
  assign rx_pin[128] = mb1_FA1_TA1_IO_116_mb1_FB1_TA2_IO_114;
  assign rx_pin[129] = mb1_FA1_TA1_IO_117_mb1_FB1_TA2_IO_115;
  assign rx_pin[130] = mb1_FA1_TA1_IO_118_mb1_FB1_TA2_IO_132;
  assign rx_pin[131] = mb1_FA1_TA1_IO_119_mb1_FB1_TA2_IO_133;
  assign rx_pin[132] = mb1_FA1_TA1_IO_120_mb1_FB1_TA2_IO_130;
  assign rx_pin[133] = mb1_FA1_TA1_IO_121_mb1_FB1_TA2_IO_131;
  assign rx_pin[134] = mb1_FA1_TA1_IO_122_mb1_FB1_TA2_IO_108;
  assign rx_pin[135] = mb1_FA1_TA1_IO_123_mb1_FB1_TA2_IO_109;
  assign rx_pin[136] = mb1_FA1_TA1_IO_124_mb1_FB1_TA2_IO_126;
  assign rx_pin[137] = mb1_FA1_TA1_IO_125_mb1_FB1_TA2_IO_127;
  assign rx_pin[138] = mb1_FA1_TA1_IO_126_mb1_FB1_TA2_IO_124;
  assign rx_pin[139] = mb1_FA1_TA1_IO_127_mb1_FB1_TA2_IO_125;
  assign rx_pin[140] = mb1_FA1_TA1_IO_130_mb1_FB1_TA2_IO_120;
  assign rx_pin[141] = mb1_FA1_TA1_IO_131_mb1_FB1_TA2_IO_121;
  assign rx_pin[142] = mb1_FA1_TA1_IO_132_mb1_FB1_TA2_IO_118;
  assign rx_pin[143] = mb1_FA1_TA1_IO_133_mb1_FB1_TA2_IO_119;
  assign rx_pin[144] = mb1_FA1_TA1_IO_134_mb1_FB1_TA2_IO_136;
  assign rx_pin[145] = mb1_FA1_TA1_IO_136_mb1_FB1_TA2_IO_134;
  assign mb1_FB1_TB0_CLKIO_N_0_mb1_FB2_BB2_CLKIO_N_7 = tx_pin[146];
  assign mb1_FB1_TB0_CLKIO_N_1_mb1_FB2_BB2_CLKIO_N_6 = tx_pin[147];
  assign mb1_FB1_TB0_CLKIO_N_2_mb1_FB2_BB2_CLKIO_N_4 = tx_pin[148];
  assign mb1_FB1_TB0_CLKIO_N_3_mb1_FB2_BB2_CLKIO_N_3 = tx_pin[149];
  assign mb1_FB1_TB0_CLKIO_N_4_mb1_FB2_BB2_CLKIO_N_2 = tx_pin[150];
  assign mb1_FB1_TB0_CLKIO_N_5_mb1_FB2_BB2_IO_010 = tx_pin[151];
  assign mb1_FB1_TB0_CLKIO_N_6_mb1_FB2_BB2_CLKIO_N_1 = tx_pin[152];
  assign mb1_FB1_TB0_CLKIO_N_7_mb1_FB2_BB2_CLKIO_N_0 = tx_pin[153];
  assign mb1_FB1_TB0_CLKIO_P_0_mb1_FB2_BB2_CLKIO_P_7 = tx_pin[154];
  assign mb1_FB1_TB0_CLKIO_P_1_mb1_FB2_BB2_CLKIO_P_6 = tx_pin[155];
  assign mb1_FB1_TB0_CLKIO_P_2_mb1_FB2_BB2_CLKIO_P_4 = tx_pin[156];
  assign mb1_FB1_TB0_CLKIO_P_3_mb1_FB2_BB2_CLKIO_P_3 = tx_pin[157];
  assign mb1_FB1_TB0_CLKIO_P_4_mb1_FB2_BB2_CLKIO_P_2 = tx_pin[158];
  assign mb1_FB1_TB0_CLKIO_P_5_mb1_FB2_BB2_IO_011 = tx_pin[159];
  assign mb1_FB1_TB0_CLKIO_P_6_mb1_FB2_BB2_CLKIO_P_1 = tx_pin[160];
  assign mb1_FB1_TB0_CLKIO_P_7_mb1_FB2_BB2_CLKIO_P_0 = tx_pin[161];
  assign mb1_FB1_TB0_IO_004_mb1_FB2_BB2_IO_006 = tx_pin[162];
  assign mb1_FB1_TB0_IO_005_mb1_FB2_BB2_IO_007 = tx_pin[163];
  assign mb1_FB1_TB0_IO_006_mb1_FB2_BB2_IO_004 = tx_pin[164];
  assign mb1_FB1_TB0_IO_007_mb1_FB2_BB2_IO_005 = tx_pin[165];
  assign mb1_FB1_TB0_IO_008_mb1_FB2_BB2_IO_022 = tx_pin[166];
  assign mb1_FB1_TB0_IO_009_mb1_FB2_BB2_IO_023 = tx_pin[167];
  assign mb1_FB1_TB0_IO_010_mb1_FB2_BB2_CLKIO_N_5 = tx_pin[168];
  assign mb1_FB1_TB0_IO_011_mb1_FB2_BB2_CLKIO_P_5 = tx_pin[169];
  assign mb1_FB1_TB0_IO_012_mb1_FB2_BB2_IO_012 = tx_pin[170];
  assign mb1_FB1_TB0_IO_013_mb1_FB2_BB2_IO_013 = tx_pin[171];
  assign mb1_FB1_TB0_IO_014_mb1_FB2_BB2_IO_016 = tx_pin[172];
  assign mb1_FB1_TB0_IO_015_mb1_FB2_BB2_IO_017 = tx_pin[173];
  assign mb1_FB1_TB0_IO_016_mb1_FB2_BB2_IO_014 = tx_pin[174];
  assign mb1_FB1_TB0_IO_017_mb1_FB2_BB2_IO_015 = tx_pin[175];
  assign mb1_FB1_TB0_IO_018_mb1_FB2_BB2_IO_032 = tx_pin[176];
  assign mb1_FB1_TB0_IO_019_mb1_FB2_BB2_IO_033 = tx_pin[177];
  assign mb1_FB1_TB0_IO_020_mb1_FB2_BB2_IO_030 = tx_pin[178];
  assign mb1_FB1_TB0_IO_021_mb1_FB2_BB2_IO_031 = tx_pin[179];
  assign mb1_FB1_TB0_IO_022_mb1_FB2_BB2_IO_008 = tx_pin[180];
  assign mb1_FB1_TB0_IO_023_mb1_FB2_BB2_IO_009 = tx_pin[181];
  assign mb1_FB1_TB0_IO_024_mb1_FB2_BB2_IO_026 = tx_pin[182];
  assign mb1_FB1_TB0_IO_025_mb1_FB2_BB2_IO_027 = tx_pin[183];
  assign mb1_FB1_TB0_IO_026_mb1_FB2_BB2_IO_024 = tx_pin[184];
  assign mb1_FB1_TB0_IO_027_mb1_FB2_BB2_IO_025 = tx_pin[185];
  assign mb1_FB1_TB0_IO_028_mb1_FB2_BB2_IO_042 = tx_pin[186];
  assign mb1_FB1_TB0_IO_029_mb1_FB2_BB2_IO_043 = tx_pin[187];
  assign mb1_FB1_TB0_IO_030_mb1_FB2_BB2_IO_020 = tx_pin[188];
  assign mb1_FB1_TB0_IO_031_mb1_FB2_BB2_IO_021 = tx_pin[189];
  assign mb1_FB1_TB0_IO_032_mb1_FB2_BB2_IO_018 = tx_pin[190];
  assign mb1_FB1_TB0_IO_033_mb1_FB2_BB2_IO_019 = tx_pin[191];
  assign mb1_FB1_TB0_IO_034_mb1_FB2_BB2_IO_036 = tx_pin[192];
  assign mb1_FB1_TB0_IO_035_mb1_FB2_BB2_IO_037 = tx_pin[193];
  assign mb1_FB1_TB0_IO_036_mb1_FB2_BB2_IO_034 = tx_pin[194];
  assign mb1_FB1_TB0_IO_037_mb1_FB2_BB2_IO_035 = tx_pin[195];
  assign mb1_FB1_TB0_IO_038_mb1_FB2_BB2_IO_052 = tx_pin[196];
  assign mb1_FB1_TB0_IO_039_mb1_FB2_BB2_IO_053 = tx_pin[197];
  assign mb1_FB1_TB0_IO_040_mb1_FB2_BB2_IO_050 = tx_pin[198];
  assign mb1_FB1_TB0_IO_041_mb1_FB2_BB2_IO_051 = tx_pin[199];
  assign mb1_FB1_TB0_IO_042_mb1_FB2_BB2_IO_028 = tx_pin[200];
  assign mb1_FB1_TB0_IO_043_mb1_FB2_BB2_IO_029 = tx_pin[201];
  assign mb1_FB1_TB0_IO_044_mb1_FB2_BB2_IO_046 = tx_pin[202];
  assign mb1_FB1_TB0_IO_045_mb1_FB2_BB2_IO_047 = tx_pin[203];
  assign mb1_FB1_TB0_IO_046_mb1_FB2_BB2_IO_044 = tx_pin[204];
  assign mb1_FB1_TB0_IO_047_mb1_FB2_BB2_IO_045 = tx_pin[205];
  assign mb1_FB1_TB0_IO_048_mb1_FB2_BB2_IO_062 = tx_pin[206];
  assign mb1_FB1_TB0_IO_049_mb1_FB2_BB2_IO_063 = tx_pin[207];
  assign mb1_FB1_TB0_IO_050_mb1_FB2_BB2_IO_040 = tx_pin[208];
  assign mb1_FB1_TB0_IO_051_mb1_FB2_BB2_IO_041 = tx_pin[209];
  assign mb1_FB1_TB0_IO_052_mb1_FB2_BB2_IO_038 = tx_pin[210];
  assign mb1_FB1_TB0_IO_053_mb1_FB2_BB2_IO_039 = tx_pin[211];
  assign mb1_FB1_TB0_IO_054_mb1_FB2_BB2_IO_056 = tx_pin[212];
  assign mb1_FB1_TB0_IO_055_mb1_FB2_BB2_IO_057 = tx_pin[213];
  assign mb1_FB1_TB0_IO_056_mb1_FB2_BB2_IO_054 = tx_pin[214];
  assign mb1_FB1_TB0_IO_057_mb1_FB2_BB2_IO_055 = tx_pin[215];
  assign mb1_FB1_TB0_IO_058_mb1_FB2_BB2_IO_072 = tx_pin[216];
  assign mb1_FB1_TB0_IO_059_mb1_FB2_BB2_IO_073 = tx_pin[217];
  assign mb1_FB1_TB0_IO_060_mb1_FB2_BB2_IO_070 = tx_pin[218];
  assign mb1_FB1_TB0_IO_061_mb1_FB2_BB2_IO_071 = tx_pin[219];
  assign mb1_FB1_TB0_IO_062_mb1_FB2_BB2_IO_048 = tx_pin[220];
  assign mb1_FB1_TB0_IO_063_mb1_FB2_BB2_IO_049 = tx_pin[221];
  assign mb1_FB1_TB0_IO_064_mb1_FB2_BB2_IO_066 = tx_pin[222];
  assign mb1_FB1_TB0_IO_065_mb1_FB2_BB2_IO_067 = tx_pin[223];
  assign mb1_FB1_TB0_IO_066_mb1_FB2_BB2_IO_064 = tx_pin[224];
  assign mb1_FB1_TB0_IO_067_mb1_FB2_BB2_IO_065 = tx_pin[225];
  assign mb1_FB1_TB0_IO_068_mb1_FB2_BB2_IO_082 = tx_pin[226];
  assign mb1_FB1_TB0_IO_069_mb1_FB2_BB2_IO_083 = tx_pin[227];
  assign mb1_FB1_TB0_IO_070_mb1_FB2_BB2_IO_060 = tx_pin[228];
  assign mb1_FB1_TB0_IO_071_mb1_FB2_BB2_IO_061 = tx_pin[229];
  assign mb1_FB1_TB0_IO_072_mb1_FB2_BB2_IO_058 = tx_pin[230];
  assign mb1_FB1_TB0_IO_073_mb1_FB2_BB2_IO_059 = tx_pin[231];
  assign mb1_FB1_TB0_IO_074_mb1_FB2_BB2_IO_076 = tx_pin[232];
  assign mb1_FB1_TB0_IO_075_mb1_FB2_BB2_IO_077 = tx_pin[233];
  assign mb1_FB1_TB0_IO_076_mb1_FB2_BB2_IO_074 = tx_pin[234];
  assign mb1_FB1_TB0_IO_077_mb1_FB2_BB2_IO_075 = tx_pin[235];
  assign mb1_FB1_TB0_IO_078_mb1_FB2_BB2_IO_092 = tx_pin[236];
  assign mb1_FB1_TB0_IO_079_mb1_FB2_BB2_IO_093 = tx_pin[237];
  assign mb1_FB1_TB0_IO_080_mb1_FB2_BB2_IO_090 = tx_pin[238];
  assign mb1_FB1_TB0_IO_081_mb1_FB2_BB2_IO_091 = tx_pin[239];
  assign mb1_FB1_TB0_IO_082_mb1_FB2_BB2_IO_068 = tx_pin[240];
  assign mb1_FB1_TB0_IO_083_mb1_FB2_BB2_IO_069 = tx_pin[241];
  assign mb1_FB1_TB0_IO_084_mb1_FB2_BB2_IO_086 = tx_pin[242];
  assign mb1_FB1_TB0_IO_085_mb1_FB2_BB2_IO_087 = tx_pin[243];
  assign mb1_FB1_TB0_IO_086_mb1_FB2_BB2_IO_084 = tx_pin[244];
  assign mb1_FB1_TB0_IO_087_mb1_FB2_BB2_IO_085 = tx_pin[245];
  assign mb1_FB1_TB0_IO_088_mb1_FB2_BB2_IO_102 = tx_pin[246];
  assign mb1_FB1_TB0_IO_089_mb1_FB2_BB2_IO_103 = tx_pin[247];
  assign mb1_FB1_TB0_IO_090_mb1_FB2_BB2_IO_080 = tx_pin[248];
  assign mb1_FB1_TB0_IO_091_mb1_FB2_BB2_IO_081 = tx_pin[249];
  assign mb1_FB1_TB0_IO_092_mb1_FB2_BB2_IO_078 = tx_pin[250];
  assign mb1_FB1_TB0_IO_093_mb1_FB2_BB2_IO_079 = tx_pin[251];
  assign mb1_FB1_TB0_IO_094_mb1_FB2_BB2_IO_096 = tx_pin[252];
  assign mb1_FB1_TB0_IO_095_mb1_FB2_BB2_IO_097 = tx_pin[253];
  assign mb1_FB1_TB0_IO_096_mb1_FB2_BB2_IO_094 = tx_pin[254];
  assign mb1_FB1_TB0_IO_097_mb1_FB2_BB2_IO_095 = tx_pin[255];
  assign mb1_FB1_TB0_IO_098_mb1_FB2_BB2_IO_112 = tx_pin[256];
  assign mb1_FB1_TB0_IO_099_mb1_FB2_BB2_IO_113 = tx_pin[257];
  assign mb1_FB1_TB0_IO_100_mb1_FB2_BB2_IO_110 = tx_pin[258];
  assign mb1_FB1_TB0_IO_101_mb1_FB2_BB2_IO_111 = tx_pin[259];
  assign mb1_FB1_TB0_IO_102_mb1_FB2_BB2_IO_088 = tx_pin[260];
  assign mb1_FB1_TB0_IO_103_mb1_FB2_BB2_IO_089 = tx_pin[261];
  assign mb1_FB1_TB0_IO_104_mb1_FB2_BB2_IO_106 = tx_pin[262];
  assign mb1_FB1_TB0_IO_105_mb1_FB2_BB2_IO_107 = tx_pin[263];
  assign mb1_FB1_TB0_IO_106_mb1_FB2_BB2_IO_104 = tx_pin[264];
  assign mb1_FB1_TB0_IO_107_mb1_FB2_BB2_IO_105 = tx_pin[265];
  assign mb1_FB1_TB0_IO_108_mb1_FB2_BB2_IO_122 = tx_pin[266];
  assign mb1_FB1_TB0_IO_109_mb1_FB2_BB2_IO_123 = tx_pin[267];
  assign mb1_FB1_TB0_IO_110_mb1_FB2_BB2_IO_100 = tx_pin[268];
  assign mb1_FB1_TB0_IO_111_mb1_FB2_BB2_IO_101 = tx_pin[269];
  assign mb1_FB1_TB0_IO_112_mb1_FB2_BB2_IO_098 = tx_pin[270];
  assign mb1_FB1_TB0_IO_113_mb1_FB2_BB2_IO_099 = tx_pin[271];
  assign mb1_FB1_TB0_IO_114_mb1_FB2_BB2_IO_116 = tx_pin[272];
  assign mb1_FB1_TB0_IO_115_mb1_FB2_BB2_IO_117 = tx_pin[273];
  assign mb1_FB1_TB0_IO_116_mb1_FB2_BB2_IO_114 = tx_pin[274];
  assign mb1_FB1_TB0_IO_117_mb1_FB2_BB2_IO_115 = tx_pin[275];
  assign mb1_FB1_TB0_IO_118_mb1_FB2_BB2_IO_132 = tx_pin[276];
  assign mb1_FB1_TB0_IO_119_mb1_FB2_BB2_IO_133 = tx_pin[277];
  assign mb1_FB1_TB0_IO_120_mb1_FB2_BB2_IO_130 = tx_pin[278];
  assign mb1_FB1_TB0_IO_121_mb1_FB2_BB2_IO_131 = tx_pin[279];
  assign mb1_FB1_TB0_IO_122_mb1_FB2_BB2_IO_108 = tx_pin[280];
  assign mb1_FB1_TB0_IO_123_mb1_FB2_BB2_IO_109 = tx_pin[281];
  assign mb1_FB1_TB0_IO_124_mb1_FB2_BB2_IO_126 = tx_pin[282];
  assign mb1_FB1_TB0_IO_125_mb1_FB2_BB2_IO_127 = tx_pin[283];
  assign mb1_FB1_TB0_IO_126_mb1_FB2_BB2_IO_124 = tx_pin[284];
  assign mb1_FB1_TB0_IO_127_mb1_FB2_BB2_IO_125 = tx_pin[285];
  assign mb1_FB1_TB0_IO_130_mb1_FB2_BB2_IO_120 = tx_pin[286];
  assign mb1_FB1_TB0_IO_131_mb1_FB2_BB2_IO_121 = tx_pin[287];
  assign mb1_FB1_TB0_IO_132_mb1_FB2_BB2_IO_118 = tx_pin[288];
  assign mb1_FB1_TB0_IO_133_mb1_FB2_BB2_IO_119 = tx_pin[289];
  assign mb1_FB1_TB0_IO_134_mb1_FB2_BB2_IO_136 = tx_pin[290];
  assign mb1_FB1_TB0_IO_136_mb1_FB2_BB2_IO_134 = tx_pin[291];
  assign mb1_FB1_TB1_CLKIO_N_0_mb1_FA2_BA1_CLKIO_N_7 = tx_pin[292];
  assign mb1_FB1_TB1_CLKIO_N_1_mb1_FA2_BA1_CLKIO_N_6 = tx_pin[293];
  assign mb1_FB1_TB1_CLKIO_N_2_mb1_FA2_BA1_CLKIO_N_4 = tx_pin[294];
  assign mb1_FB1_TB1_CLKIO_N_3_mb1_FA2_BA1_CLKIO_N_3 = tx_pin[295];
  assign mb1_FB1_TB1_CLKIO_N_4_mb1_FA2_BA1_CLKIO_N_2 = tx_pin[296];
  assign mb1_FB1_TB1_CLKIO_N_5_mb1_FA2_BA1_IO_010 = tx_pin[297];
  assign mb1_FB1_TB1_CLKIO_N_6_mb1_FA2_BA1_CLKIO_N_1 = tx_pin[298];
  assign mb1_FB1_TB1_CLKIO_N_7_mb1_FA2_BA1_CLKIO_N_0 = tx_pin[299];
  assign mb1_FB1_TB1_CLKIO_P_0_mb1_FA2_BA1_CLKIO_P_7 = tx_pin[300];
  assign mb1_FB1_TB1_CLKIO_P_1_mb1_FA2_BA1_CLKIO_P_6 = tx_pin[301];
  assign mb1_FB1_TB1_CLKIO_P_2_mb1_FA2_BA1_CLKIO_P_4 = tx_pin[302];
  assign mb1_FB1_TB1_CLKIO_P_3_mb1_FA2_BA1_CLKIO_P_3 = tx_pin[303];
  assign mb1_FB1_TB1_CLKIO_P_4_mb1_FA2_BA1_CLKIO_P_2 = tx_pin[304];
  assign mb1_FB1_TB1_CLKIO_P_5_mb1_FA2_BA1_IO_011 = tx_pin[305];
  assign mb1_FB1_TB1_CLKIO_P_6_mb1_FA2_BA1_CLKIO_P_1 = tx_pin[306];
  assign mb1_FB1_TB1_CLKIO_P_7_mb1_FA2_BA1_CLKIO_P_0 = tx_pin[307];
  assign mb1_FB1_TB1_IO_004_mb1_FA2_BA1_IO_006 = tx_pin[308];
  assign mb1_FB1_TB1_IO_005_mb1_FA2_BA1_IO_007 = tx_pin[309];
  assign mb1_FB1_TB1_IO_006_mb1_FA2_BA1_IO_004 = tx_pin[310];
  assign mb1_FB1_TB1_IO_007_mb1_FA2_BA1_IO_005 = tx_pin[311];
  assign mb1_FB1_TB1_IO_008_mb1_FA2_BA1_IO_022 = tx_pin[312];
  assign mb1_FB1_TB1_IO_009_mb1_FA2_BA1_IO_023 = tx_pin[313];
  assign mb1_FB1_TB1_IO_010_mb1_FA2_BA1_CLKIO_N_5 = tx_pin[314];
  assign mb1_FB1_TB1_IO_011_mb1_FA2_BA1_CLKIO_P_5 = tx_pin[315];
  assign mb1_FB1_TB1_IO_012_mb1_FA2_BA1_IO_012 = tx_pin[316];
  assign mb1_FB1_TB1_IO_013_mb1_FA2_BA1_IO_013 = tx_pin[317];
  assign mb1_FB1_TB1_IO_014_mb1_FA2_BA1_IO_016 = tx_pin[318];
  assign mb1_FB1_TB1_IO_015_mb1_FA2_BA1_IO_017 = tx_pin[319];
  assign mb1_FB1_TB1_IO_016_mb1_FA2_BA1_IO_014 = tx_pin[320];
  assign mb1_FB1_TB1_IO_017_mb1_FA2_BA1_IO_015 = tx_pin[321];
  assign mb1_FB1_TB1_IO_018_mb1_FA2_BA1_IO_032 = tx_pin[322];
  assign mb1_FB1_TB1_IO_019_mb1_FA2_BA1_IO_033 = tx_pin[323];
  assign mb1_FB1_TB1_IO_020_mb1_FA2_BA1_IO_030 = tx_pin[324];
  assign mb1_FB1_TB1_IO_021_mb1_FA2_BA1_IO_031 = tx_pin[325];
  assign mb1_FB1_TB1_IO_022_mb1_FA2_BA1_IO_008 = tx_pin[326];
  assign mb1_FB1_TB1_IO_023_mb1_FA2_BA1_IO_009 = tx_pin[327];
  assign mb1_FB1_TB1_IO_024_mb1_FA2_BA1_IO_026 = tx_pin[328];
  assign mb1_FB1_TB1_IO_025_mb1_FA2_BA1_IO_027 = tx_pin[329];
  assign mb1_FB1_TB1_IO_026_mb1_FA2_BA1_IO_024 = tx_pin[330];
  assign mb1_FB1_TB1_IO_027_mb1_FA2_BA1_IO_025 = tx_pin[331];
  assign mb1_FB1_TB1_IO_028_mb1_FA2_BA1_IO_042 = tx_pin[332];
  assign mb1_FB1_TB1_IO_029_mb1_FA2_BA1_IO_043 = tx_pin[333];
  assign mb1_FB1_TB1_IO_030_mb1_FA2_BA1_IO_020 = tx_pin[334];
  assign mb1_FB1_TB1_IO_031_mb1_FA2_BA1_IO_021 = tx_pin[335];
  assign mb1_FB1_TB1_IO_032_mb1_FA2_BA1_IO_018 = tx_pin[336];
  assign mb1_FB1_TB1_IO_033_mb1_FA2_BA1_IO_019 = tx_pin[337];
  assign mb1_FB1_TB1_IO_034_mb1_FA2_BA1_IO_036 = tx_pin[338];
  assign mb1_FB1_TB1_IO_035_mb1_FA2_BA1_IO_037 = tx_pin[339];
  assign mb1_FB1_TB1_IO_036_mb1_FA2_BA1_IO_034 = tx_pin[340];
  assign mb1_FB1_TB1_IO_037_mb1_FA2_BA1_IO_035 = tx_pin[341];
  assign mb1_FB1_TB1_IO_038_mb1_FA2_BA1_IO_052 = tx_pin[342];
  assign mb1_FB1_TB1_IO_039_mb1_FA2_BA1_IO_053 = tx_pin[343];
  assign mb1_FB1_TB1_IO_040_mb1_FA2_BA1_IO_050 = tx_pin[344];
  assign mb1_FB1_TB1_IO_041_mb1_FA2_BA1_IO_051 = tx_pin[345];
  assign mb1_FB1_TB1_IO_042_mb1_FA2_BA1_IO_028 = tx_pin[346];
  assign mb1_FB1_TB1_IO_043_mb1_FA2_BA1_IO_029 = tx_pin[347];
  assign mb1_FB1_TB1_IO_044_mb1_FA2_BA1_IO_046 = tx_pin[348];
  assign mb1_FB1_TB1_IO_045_mb1_FA2_BA1_IO_047 = tx_pin[349];
  assign mb1_FB1_TB1_IO_046_mb1_FA2_BA1_IO_044 = tx_pin[350];
  assign mb1_FB1_TB1_IO_047_mb1_FA2_BA1_IO_045 = tx_pin[351];
  assign mb1_FB1_TB1_IO_048_mb1_FA2_BA1_IO_062 = tx_pin[352];
  assign mb1_FB1_TB1_IO_049_mb1_FA2_BA1_IO_063 = tx_pin[353];
  assign mb1_FB1_TB1_IO_050_mb1_FA2_BA1_IO_040 = tx_pin[354];
  assign mb1_FB1_TB1_IO_051_mb1_FA2_BA1_IO_041 = tx_pin[355];
  assign mb1_FB1_TB1_IO_052_mb1_FA2_BA1_IO_038 = tx_pin[356];
  assign mb1_FB1_TB1_IO_053_mb1_FA2_BA1_IO_039 = tx_pin[357];
  assign mb1_FB1_TB1_IO_054_mb1_FA2_BA1_IO_056 = tx_pin[358];
  assign mb1_FB1_TB1_IO_055_mb1_FA2_BA1_IO_057 = tx_pin[359];
  assign mb1_FB1_TB1_IO_056_mb1_FA2_BA1_IO_054 = tx_pin[360];
  assign mb1_FB1_TB1_IO_057_mb1_FA2_BA1_IO_055 = tx_pin[361];
  assign mb1_FB1_TB1_IO_058_mb1_FA2_BA1_IO_072 = tx_pin[362];
  assign mb1_FB1_TB1_IO_059_mb1_FA2_BA1_IO_073 = tx_pin[363];
  assign mb1_FB1_TB1_IO_060_mb1_FA2_BA1_IO_070 = tx_pin[364];
  assign mb1_FB1_TB1_IO_061_mb1_FA2_BA1_IO_071 = tx_pin[365];
  assign mb1_FB1_TB1_IO_062_mb1_FA2_BA1_IO_048 = tx_pin[366];
  assign mb1_FB1_TB1_IO_063_mb1_FA2_BA1_IO_049 = tx_pin[367];
  assign mb1_FB1_TB1_IO_064_mb1_FA2_BA1_IO_066 = tx_pin[368];
  assign mb1_FB1_TB1_IO_065_mb1_FA2_BA1_IO_067 = tx_pin[369];
  assign mb1_FB1_TB1_IO_066_mb1_FA2_BA1_IO_064 = tx_pin[370];
  assign mb1_FB1_TB1_IO_067_mb1_FA2_BA1_IO_065 = tx_pin[371];
  assign mb1_FB1_TB1_IO_068_mb1_FA2_BA1_IO_082 = tx_pin[372];
  assign mb1_FB1_TB1_IO_069_mb1_FA2_BA1_IO_083 = tx_pin[373];
  assign mb1_FB1_TB1_IO_070_mb1_FA2_BA1_IO_060 = tx_pin[374];
  assign mb1_FB1_TB1_IO_071_mb1_FA2_BA1_IO_061 = tx_pin[375];
  assign mb1_FB1_TB1_IO_072_mb1_FA2_BA1_IO_058 = tx_pin[376];
  assign mb1_FB1_TB1_IO_073_mb1_FA2_BA1_IO_059 = tx_pin[377];
  assign mb1_FB1_TB1_IO_074_mb1_FA2_BA1_IO_076 = tx_pin[378];
  assign mb1_FB1_TB1_IO_075_mb1_FA2_BA1_IO_077 = tx_pin[379];
  assign mb1_FB1_TB1_IO_076_mb1_FA2_BA1_IO_074 = tx_pin[380];
  assign mb1_FB1_TB1_IO_077_mb1_FA2_BA1_IO_075 = tx_pin[381];
  assign mb1_FB1_TB1_IO_078_mb1_FA2_BA1_IO_092 = tx_pin[382];
  assign mb1_FB1_TB1_IO_079_mb1_FA2_BA1_IO_093 = tx_pin[383];
  assign mb1_FB1_TB1_IO_080_mb1_FA2_BA1_IO_090 = tx_pin[384];
  assign mb1_FB1_TB1_IO_081_mb1_FA2_BA1_IO_091 = tx_pin[385];
  assign mb1_FB1_TB1_IO_082_mb1_FA2_BA1_IO_068 = tx_pin[386];
  assign mb1_FB1_TB1_IO_083_mb1_FA2_BA1_IO_069 = tx_pin[387];
  assign mb1_FB1_TB1_IO_084_mb1_FA2_BA1_IO_086 = tx_pin[388];
  assign mb1_FB1_TB1_IO_085_mb1_FA2_BA1_IO_087 = tx_pin[389];
  assign mb1_FB1_TB1_IO_086_mb1_FA2_BA1_IO_084 = tx_pin[390];
  assign mb1_FB1_TB1_IO_087_mb1_FA2_BA1_IO_085 = tx_pin[391];
  assign mb1_FB1_TB1_IO_088_mb1_FA2_BA1_IO_102 = tx_pin[392];
  assign mb1_FB1_TB1_IO_089_mb1_FA2_BA1_IO_103 = tx_pin[393];
  assign mb1_FB1_TB1_IO_090_mb1_FA2_BA1_IO_080 = tx_pin[394];
  assign mb1_FB1_TB1_IO_091_mb1_FA2_BA1_IO_081 = tx_pin[395];
  assign mb1_FB1_TB1_IO_092_mb1_FA2_BA1_IO_078 = tx_pin[396];
  assign mb1_FB1_TB1_IO_093_mb1_FA2_BA1_IO_079 = tx_pin[397];
  assign mb1_FB1_TB1_IO_094_mb1_FA2_BA1_IO_096 = tx_pin[398];
  assign mb1_FB1_TB1_IO_095_mb1_FA2_BA1_IO_097 = tx_pin[399];
  assign mb1_FB1_TB1_IO_096_mb1_FA2_BA1_IO_094 = tx_pin[400];
  assign mb1_FB1_TB1_IO_097_mb1_FA2_BA1_IO_095 = tx_pin[401];
  assign mb1_FB1_TB1_IO_098_mb1_FA2_BA1_IO_112 = tx_pin[402];
  assign mb1_FB1_TB1_IO_099_mb1_FA2_BA1_IO_113 = tx_pin[403];
  assign mb1_FB1_TB1_IO_100_mb1_FA2_BA1_IO_110 = tx_pin[404];
  assign mb1_FB1_TB1_IO_101_mb1_FA2_BA1_IO_111 = tx_pin[405];
  assign mb1_FB1_TB1_IO_102_mb1_FA2_BA1_IO_088 = tx_pin[406];
  assign mb1_FB1_TB1_IO_103_mb1_FA2_BA1_IO_089 = tx_pin[407];
  assign mb1_FB1_TB1_IO_104_mb1_FA2_BA1_IO_106 = tx_pin[408];
  assign mb1_FB1_TB1_IO_105_mb1_FA2_BA1_IO_107 = tx_pin[409];
  assign mb1_FB1_TB1_IO_106_mb1_FA2_BA1_IO_104 = tx_pin[410];
  assign mb1_FB1_TB1_IO_107_mb1_FA2_BA1_IO_105 = tx_pin[411];
  assign mb1_FB1_TB1_IO_108_mb1_FA2_BA1_IO_122 = tx_pin[412];
  assign mb1_FB1_TB1_IO_109_mb1_FA2_BA1_IO_123 = tx_pin[413];
  assign mb1_FB1_TB1_IO_110_mb1_FA2_BA1_IO_100 = tx_pin[414];
  assign mb1_FB1_TB1_IO_111_mb1_FA2_BA1_IO_101 = tx_pin[415];
  assign mb1_FB1_TB1_IO_112_mb1_FA2_BA1_IO_098 = tx_pin[416];
  assign mb1_FB1_TB1_IO_113_mb1_FA2_BA1_IO_099 = tx_pin[417];
  assign mb1_FB1_TB1_IO_114_mb1_FA2_BA1_IO_116 = tx_pin[418];
  assign mb1_FB1_TB1_IO_115_mb1_FA2_BA1_IO_117 = tx_pin[419];
  assign mb1_FB1_TB1_IO_116_mb1_FA2_BA1_IO_114 = tx_pin[420];
  assign mb1_FB1_TB1_IO_117_mb1_FA2_BA1_IO_115 = tx_pin[421];
  assign mb1_FB1_TB1_IO_118_mb1_FA2_BA1_IO_132 = tx_pin[422];
  assign mb1_FB1_TB1_IO_119_mb1_FA2_BA1_IO_133 = tx_pin[423];
  assign mb1_FB1_TB1_IO_120_mb1_FA2_BA1_IO_130 = tx_pin[424];
  assign mb1_FB1_TB1_IO_121_mb1_FA2_BA1_IO_131 = tx_pin[425];
  assign mb1_FB1_TB1_IO_122_mb1_FA2_BA1_IO_108 = tx_pin[426];
  assign mb1_FB1_TB1_IO_123_mb1_FA2_BA1_IO_109 = tx_pin[427];
  assign mb1_FB1_TB1_IO_124_mb1_FA2_BA1_IO_126 = tx_pin[428];
  assign mb1_FB1_TB1_IO_125_mb1_FA2_BA1_IO_127 = tx_pin[429];
  assign mb1_FB1_TB1_IO_126_mb1_FA2_BA1_IO_124 = tx_pin[430];
  assign mb1_FB1_TB1_IO_127_mb1_FA2_BA1_IO_125 = tx_pin[431];
  assign mb1_FB1_TB1_IO_130_mb1_FA2_BA1_IO_120 = tx_pin[432];
  assign mb1_FB1_TB1_IO_131_mb1_FA2_BA1_IO_121 = tx_pin[433];
  assign mb1_FB1_TB1_IO_132_mb1_FA2_BA1_IO_118 = tx_pin[434];
  assign mb1_FB1_TB1_IO_133_mb1_FA2_BA1_IO_119 = tx_pin[435];
  assign mb1_FB1_TB1_IO_134_mb1_FA2_BA1_IO_136 = tx_pin[436];
  assign mb1_FB1_TB1_IO_136_mb1_FA2_BA1_IO_134 = tx_pin[437];
  assign rx_pin[146] = mb1_FA1_TB0_CLKIO_N_0_mb1_FB1_TB2_CLKIO_N_7;
  assign rx_pin[147] = mb1_FA1_TB0_CLKIO_N_1_mb1_FB1_TB2_CLKIO_N_6;
  assign rx_pin[148] = mb1_FA1_TB0_CLKIO_N_2_mb1_FB1_TB2_CLKIO_N_4;
  assign rx_pin[149] = mb1_FA1_TB0_CLKIO_N_3_mb1_FB1_TB2_CLKIO_N_3;
  assign rx_pin[150] = mb1_FA1_TB0_CLKIO_N_4_mb1_FB1_TB2_CLKIO_N_2;
  assign rx_pin[151] = mb1_FA1_TB0_CLKIO_N_5_mb1_FB1_TB2_IO_010;
  assign rx_pin[152] = mb1_FA1_TB0_CLKIO_N_6_mb1_FB1_TB2_CLKIO_N_1;
  assign rx_pin[153] = mb1_FA1_TB0_CLKIO_N_7_mb1_FB1_TB2_CLKIO_N_0;
  assign rx_pin[154] = mb1_FA1_TB0_CLKIO_P_0_mb1_FB1_TB2_CLKIO_P_7;
  assign rx_pin[155] = mb1_FA1_TB0_CLKIO_P_1_mb1_FB1_TB2_CLKIO_P_6;
  assign rx_pin[156] = mb1_FA1_TB0_CLKIO_P_2_mb1_FB1_TB2_CLKIO_P_4;
  assign rx_pin[157] = mb1_FA1_TB0_CLKIO_P_3_mb1_FB1_TB2_CLKIO_P_3;
  assign rx_pin[158] = mb1_FA1_TB0_CLKIO_P_4_mb1_FB1_TB2_CLKIO_P_2;
  assign rx_pin[159] = mb1_FA1_TB0_CLKIO_P_5_mb1_FB1_TB2_IO_011;
  assign rx_pin[160] = mb1_FA1_TB0_CLKIO_P_6_mb1_FB1_TB2_CLKIO_P_1;
  assign rx_pin[161] = mb1_FA1_TB0_CLKIO_P_7_mb1_FB1_TB2_CLKIO_P_0;
  assign rx_pin[162] = mb1_FA1_TB0_IO_004_mb1_FB1_TB2_IO_006;
  assign rx_pin[163] = mb1_FA1_TB0_IO_005_mb1_FB1_TB2_IO_007;
  assign rx_pin[164] = mb1_FA1_TB0_IO_006_mb1_FB1_TB2_IO_004;
  assign rx_pin[165] = mb1_FA1_TB0_IO_007_mb1_FB1_TB2_IO_005;
  assign rx_pin[166] = mb1_FA1_TB0_IO_008_mb1_FB1_TB2_IO_022;
  assign rx_pin[167] = mb1_FA1_TB0_IO_009_mb1_FB1_TB2_IO_023;
  assign rx_pin[168] = mb1_FA1_TB0_IO_010_mb1_FB1_TB2_CLKIO_N_5;
  assign rx_pin[169] = mb1_FA1_TB0_IO_011_mb1_FB1_TB2_CLKIO_P_5;
  assign rx_pin[170] = mb1_FA1_TB0_IO_012_mb1_FB1_TB2_IO_012;
  assign rx_pin[171] = mb1_FA1_TB0_IO_013_mb1_FB1_TB2_IO_013;
  assign rx_pin[172] = mb1_FA1_TB0_IO_014_mb1_FB1_TB2_IO_016;
  assign rx_pin[173] = mb1_FA1_TB0_IO_015_mb1_FB1_TB2_IO_017;
  assign rx_pin[174] = mb1_FA1_TB0_IO_016_mb1_FB1_TB2_IO_014;
  assign rx_pin[175] = mb1_FA1_TB0_IO_017_mb1_FB1_TB2_IO_015;
  assign rx_pin[176] = mb1_FA1_TB0_IO_018_mb1_FB1_TB2_IO_032;
  assign rx_pin[177] = mb1_FA1_TB0_IO_019_mb1_FB1_TB2_IO_033;
  assign rx_pin[178] = mb1_FA1_TB0_IO_020_mb1_FB1_TB2_IO_030;
  assign rx_pin[179] = mb1_FA1_TB0_IO_021_mb1_FB1_TB2_IO_031;
  assign rx_pin[180] = mb1_FA1_TB0_IO_022_mb1_FB1_TB2_IO_008;
  assign rx_pin[181] = mb1_FA1_TB0_IO_023_mb1_FB1_TB2_IO_009;
  assign rx_pin[182] = mb1_FA1_TB0_IO_024_mb1_FB1_TB2_IO_026;
  assign rx_pin[183] = mb1_FA1_TB0_IO_025_mb1_FB1_TB2_IO_027;
  assign rx_pin[184] = mb1_FA1_TB0_IO_026_mb1_FB1_TB2_IO_024;
  assign rx_pin[185] = mb1_FA1_TB0_IO_027_mb1_FB1_TB2_IO_025;
  assign rx_pin[186] = mb1_FA1_TB0_IO_028_mb1_FB1_TB2_IO_042;
  assign rx_pin[187] = mb1_FA1_TB0_IO_029_mb1_FB1_TB2_IO_043;
  assign rx_pin[188] = mb1_FA1_TB0_IO_030_mb1_FB1_TB2_IO_020;
  assign rx_pin[189] = mb1_FA1_TB0_IO_031_mb1_FB1_TB2_IO_021;
  assign rx_pin[190] = mb1_FA1_TB0_IO_032_mb1_FB1_TB2_IO_018;
  assign rx_pin[191] = mb1_FA1_TB0_IO_033_mb1_FB1_TB2_IO_019;
  assign rx_pin[192] = mb1_FA1_TB0_IO_034_mb1_FB1_TB2_IO_036;
  assign rx_pin[193] = mb1_FA1_TB0_IO_035_mb1_FB1_TB2_IO_037;
  assign rx_pin[194] = mb1_FA1_TB0_IO_036_mb1_FB1_TB2_IO_034;
  assign rx_pin[195] = mb1_FA1_TB0_IO_037_mb1_FB1_TB2_IO_035;
  assign rx_pin[196] = mb1_FA1_TB0_IO_038_mb1_FB1_TB2_IO_052;
  assign rx_pin[197] = mb1_FA1_TB0_IO_039_mb1_FB1_TB2_IO_053;
  assign rx_pin[198] = mb1_FA1_TB0_IO_040_mb1_FB1_TB2_IO_050;
  assign rx_pin[199] = mb1_FA1_TB0_IO_041_mb1_FB1_TB2_IO_051;
  assign rx_pin[200] = mb1_FA1_TB0_IO_042_mb1_FB1_TB2_IO_028;
  assign rx_pin[201] = mb1_FA1_TB0_IO_043_mb1_FB1_TB2_IO_029;
  assign rx_pin[202] = mb1_FA1_TB0_IO_044_mb1_FB1_TB2_IO_046;
  assign rx_pin[203] = mb1_FA1_TB0_IO_045_mb1_FB1_TB2_IO_047;
  assign rx_pin[204] = mb1_FA1_TB0_IO_046_mb1_FB1_TB2_IO_044;
  assign rx_pin[205] = mb1_FA1_TB0_IO_047_mb1_FB1_TB2_IO_045;
  assign rx_pin[206] = mb1_FA1_TB0_IO_048_mb1_FB1_TB2_IO_062;
  assign rx_pin[207] = mb1_FA1_TB0_IO_049_mb1_FB1_TB2_IO_063;
  assign rx_pin[208] = mb1_FA1_TB0_IO_050_mb1_FB1_TB2_IO_040;
  assign rx_pin[209] = mb1_FA1_TB0_IO_051_mb1_FB1_TB2_IO_041;
  assign rx_pin[210] = mb1_FA1_TB0_IO_052_mb1_FB1_TB2_IO_038;
  assign rx_pin[211] = mb1_FA1_TB0_IO_053_mb1_FB1_TB2_IO_039;
  assign rx_pin[212] = mb1_FA1_TB0_IO_054_mb1_FB1_TB2_IO_056;
  assign rx_pin[213] = mb1_FA1_TB0_IO_055_mb1_FB1_TB2_IO_057;
  assign rx_pin[214] = mb1_FA1_TB0_IO_056_mb1_FB1_TB2_IO_054;
  assign rx_pin[215] = mb1_FA1_TB0_IO_057_mb1_FB1_TB2_IO_055;
  assign rx_pin[216] = mb1_FA1_TB0_IO_058_mb1_FB1_TB2_IO_072;
  assign rx_pin[217] = mb1_FA1_TB0_IO_059_mb1_FB1_TB2_IO_073;
  assign rx_pin[218] = mb1_FA1_TB0_IO_060_mb1_FB1_TB2_IO_070;
  assign rx_pin[219] = mb1_FA1_TB0_IO_061_mb1_FB1_TB2_IO_071;
  assign rx_pin[220] = mb1_FA1_TB0_IO_062_mb1_FB1_TB2_IO_048;
  assign rx_pin[221] = mb1_FA1_TB0_IO_063_mb1_FB1_TB2_IO_049;
  assign rx_pin[222] = mb1_FA1_TB0_IO_064_mb1_FB1_TB2_IO_066;
  assign rx_pin[223] = mb1_FA1_TB0_IO_065_mb1_FB1_TB2_IO_067;
  assign rx_pin[224] = mb1_FA1_TB0_IO_066_mb1_FB1_TB2_IO_064;
  assign rx_pin[225] = mb1_FA1_TB0_IO_067_mb1_FB1_TB2_IO_065;
  assign rx_pin[226] = mb1_FA1_TB0_IO_068_mb1_FB1_TB2_IO_082;
  assign rx_pin[227] = mb1_FA1_TB0_IO_069_mb1_FB1_TB2_IO_083;
  assign rx_pin[228] = mb1_FA1_TB0_IO_070_mb1_FB1_TB2_IO_060;
  assign rx_pin[229] = mb1_FA1_TB0_IO_071_mb1_FB1_TB2_IO_061;
  assign rx_pin[230] = mb1_FA1_TB0_IO_072_mb1_FB1_TB2_IO_058;
  assign rx_pin[231] = mb1_FA1_TB0_IO_073_mb1_FB1_TB2_IO_059;
  assign rx_pin[232] = mb1_FA1_TB0_IO_074_mb1_FB1_TB2_IO_076;
  assign rx_pin[233] = mb1_FA1_TB0_IO_075_mb1_FB1_TB2_IO_077;
  assign rx_pin[234] = mb1_FA1_TB0_IO_076_mb1_FB1_TB2_IO_074;
  assign rx_pin[235] = mb1_FA1_TB0_IO_077_mb1_FB1_TB2_IO_075;
  assign rx_pin[236] = mb1_FA1_TB0_IO_078_mb1_FB1_TB2_IO_092;
  assign rx_pin[237] = mb1_FA1_TB0_IO_079_mb1_FB1_TB2_IO_093;
  assign rx_pin[238] = mb1_FA1_TB0_IO_080_mb1_FB1_TB2_IO_090;
  assign rx_pin[239] = mb1_FA1_TB0_IO_081_mb1_FB1_TB2_IO_091;
  assign rx_pin[240] = mb1_FA1_TB0_IO_082_mb1_FB1_TB2_IO_068;
  assign rx_pin[241] = mb1_FA1_TB0_IO_083_mb1_FB1_TB2_IO_069;
  assign rx_pin[242] = mb1_FA1_TB0_IO_084_mb1_FB1_TB2_IO_086;
  assign rx_pin[243] = mb1_FA1_TB0_IO_085_mb1_FB1_TB2_IO_087;
  assign rx_pin[244] = mb1_FA1_TB0_IO_086_mb1_FB1_TB2_IO_084;
  assign rx_pin[245] = mb1_FA1_TB0_IO_087_mb1_FB1_TB2_IO_085;
  assign rx_pin[246] = mb1_FA1_TB0_IO_088_mb1_FB1_TB2_IO_102;
  assign rx_pin[247] = mb1_FA1_TB0_IO_089_mb1_FB1_TB2_IO_103;
  assign rx_pin[248] = mb1_FA1_TB0_IO_090_mb1_FB1_TB2_IO_080;
  assign rx_pin[249] = mb1_FA1_TB0_IO_091_mb1_FB1_TB2_IO_081;
  assign rx_pin[250] = mb1_FA1_TB0_IO_092_mb1_FB1_TB2_IO_078;
  assign rx_pin[251] = mb1_FA1_TB0_IO_093_mb1_FB1_TB2_IO_079;
  assign rx_pin[252] = mb1_FA1_TB0_IO_094_mb1_FB1_TB2_IO_096;
  assign rx_pin[253] = mb1_FA1_TB0_IO_095_mb1_FB1_TB2_IO_097;
  assign rx_pin[254] = mb1_FA1_TB0_IO_096_mb1_FB1_TB2_IO_094;
  assign rx_pin[255] = mb1_FA1_TB0_IO_097_mb1_FB1_TB2_IO_095;
  assign rx_pin[256] = mb1_FA1_TB0_IO_098_mb1_FB1_TB2_IO_112;
  assign rx_pin[257] = mb1_FA1_TB0_IO_099_mb1_FB1_TB2_IO_113;
  assign rx_pin[258] = mb1_FA1_TB0_IO_100_mb1_FB1_TB2_IO_110;
  assign rx_pin[259] = mb1_FA1_TB0_IO_101_mb1_FB1_TB2_IO_111;
  assign rx_pin[260] = mb1_FA1_TB0_IO_102_mb1_FB1_TB2_IO_088;
  assign rx_pin[261] = mb1_FA1_TB0_IO_103_mb1_FB1_TB2_IO_089;
  assign rx_pin[262] = mb1_FA1_TB0_IO_104_mb1_FB1_TB2_IO_106;
  assign rx_pin[263] = mb1_FA1_TB0_IO_105_mb1_FB1_TB2_IO_107;
  assign rx_pin[264] = mb1_FA1_TB0_IO_106_mb1_FB1_TB2_IO_104;
  assign rx_pin[265] = mb1_FA1_TB0_IO_107_mb1_FB1_TB2_IO_105;
  assign rx_pin[266] = mb1_FA1_TB0_IO_108_mb1_FB1_TB2_IO_122;
  assign rx_pin[267] = mb1_FA1_TB0_IO_109_mb1_FB1_TB2_IO_123;
  assign rx_pin[268] = mb1_FA1_TB0_IO_110_mb1_FB1_TB2_IO_100;
  assign rx_pin[269] = mb1_FA1_TB0_IO_111_mb1_FB1_TB2_IO_101;
  assign rx_pin[270] = mb1_FA1_TB0_IO_112_mb1_FB1_TB2_IO_098;
  assign rx_pin[271] = mb1_FA1_TB0_IO_113_mb1_FB1_TB2_IO_099;
  assign rx_pin[272] = mb1_FA1_TB0_IO_114_mb1_FB1_TB2_IO_116;
  assign rx_pin[273] = mb1_FA1_TB0_IO_115_mb1_FB1_TB2_IO_117;
  assign rx_pin[274] = mb1_FA1_TB0_IO_116_mb1_FB1_TB2_IO_114;
  assign rx_pin[275] = mb1_FA1_TB0_IO_117_mb1_FB1_TB2_IO_115;
  assign rx_pin[276] = mb1_FA1_TB0_IO_118_mb1_FB1_TB2_IO_132;
  assign rx_pin[277] = mb1_FA1_TB0_IO_119_mb1_FB1_TB2_IO_133;
  assign rx_pin[278] = mb1_FA1_TB0_IO_120_mb1_FB1_TB2_IO_130;
  assign rx_pin[279] = mb1_FA1_TB0_IO_121_mb1_FB1_TB2_IO_131;
  assign rx_pin[280] = mb1_FA1_TB0_IO_122_mb1_FB1_TB2_IO_108;
  assign rx_pin[281] = mb1_FA1_TB0_IO_123_mb1_FB1_TB2_IO_109;
  assign rx_pin[282] = mb1_FA1_TB0_IO_124_mb1_FB1_TB2_IO_126;
  assign rx_pin[283] = mb1_FA1_TB0_IO_125_mb1_FB1_TB2_IO_127;
  assign rx_pin[284] = mb1_FA1_TB0_IO_126_mb1_FB1_TB2_IO_124;
  assign rx_pin[285] = mb1_FA1_TB0_IO_127_mb1_FB1_TB2_IO_125;
  assign rx_pin[286] = mb1_FA1_TB0_IO_130_mb1_FB1_TB2_IO_120;
  assign rx_pin[287] = mb1_FA1_TB0_IO_131_mb1_FB1_TB2_IO_121;
  assign rx_pin[288] = mb1_FA1_TB0_IO_132_mb1_FB1_TB2_IO_118;
  assign rx_pin[289] = mb1_FA1_TB0_IO_133_mb1_FB1_TB2_IO_119;
  assign rx_pin[290] = mb1_FA1_TB0_IO_134_mb1_FB1_TB2_IO_136;
  assign rx_pin[291] = mb1_FA1_TB0_IO_136_mb1_FB1_TB2_IO_134;
  assign mb1_FB1_BA0_CLKIO_N_0_mb1_FA2_TB1_CLKIO_N_7 = tx_pin[438];
  assign mb1_FB1_BA0_CLKIO_N_1_mb1_FA2_TB1_CLKIO_N_6 = tx_pin[439];
  assign mb1_FB1_BA0_CLKIO_N_2_mb1_FA2_TB1_CLKIO_N_4 = tx_pin[440];
  assign mb1_FB1_BA0_CLKIO_N_3_mb1_FA2_TB1_CLKIO_N_3 = tx_pin[441];
  assign mb1_FB1_BA0_CLKIO_N_4_mb1_FA2_TB1_CLKIO_N_2 = tx_pin[442];
  assign mb1_FB1_BA0_CLKIO_N_5_mb1_FA2_TB1_IO_010 = tx_pin[443];
  assign mb1_FB1_BA0_CLKIO_N_6_mb1_FA2_TB1_CLKIO_N_1 = tx_pin[444];
  assign mb1_FB1_BA0_CLKIO_N_7_mb1_FA2_TB1_CLKIO_N_0 = tx_pin[445];
  assign mb1_FB1_BA0_CLKIO_P_0_mb1_FA2_TB1_CLKIO_P_7 = tx_pin[446];
  assign mb1_FB1_BA0_CLKIO_P_1_mb1_FA2_TB1_CLKIO_P_6 = tx_pin[447];
  assign mb1_FB1_BA0_CLKIO_P_2_mb1_FA2_TB1_CLKIO_P_4 = tx_pin[448];
  assign mb1_FB1_BA0_CLKIO_P_3_mb1_FA2_TB1_CLKIO_P_3 = tx_pin[449];
  assign mb1_FB1_BA0_CLKIO_P_4_mb1_FA2_TB1_CLKIO_P_2 = tx_pin[450];
  assign mb1_FB1_BA0_CLKIO_P_5_mb1_FA2_TB1_IO_011 = tx_pin[451];
  assign mb1_FB1_BA0_CLKIO_P_6_mb1_FA2_TB1_CLKIO_P_1 = tx_pin[452];
  assign mb1_FB1_BA0_CLKIO_P_7_mb1_FA2_TB1_CLKIO_P_0 = tx_pin[453];
  assign mb1_FB1_BA0_IO_004_mb1_FA2_TB1_IO_006 = tx_pin[454];
  assign mb1_FB1_BA0_IO_005_mb1_FA2_TB1_IO_007 = tx_pin[455];
  assign mb1_FB1_BA0_IO_006_mb1_FA2_TB1_IO_004 = tx_pin[456];
  assign mb1_FB1_BA0_IO_007_mb1_FA2_TB1_IO_005 = tx_pin[457];
  assign mb1_FB1_BA0_IO_008_mb1_FA2_TB1_IO_022 = tx_pin[458];
  assign mb1_FB1_BA0_IO_009_mb1_FA2_TB1_IO_023 = tx_pin[459];
  assign mb1_FB1_BA0_IO_010_mb1_FA2_TB1_CLKIO_N_5 = tx_pin[460];
  assign mb1_FB1_BA0_IO_011_mb1_FA2_TB1_CLKIO_P_5 = tx_pin[461];
  assign mb1_FB1_BA0_IO_012_mb1_FA2_TB1_IO_012 = tx_pin[462];
  assign mb1_FB1_BA0_IO_013_mb1_FA2_TB1_IO_013 = tx_pin[463];
  assign mb1_FB1_BA0_IO_014_mb1_FA2_TB1_IO_016 = tx_pin[464];
  assign mb1_FB1_BA0_IO_015_mb1_FA2_TB1_IO_017 = tx_pin[465];
  assign mb1_FB1_BA0_IO_016_mb1_FA2_TB1_IO_014 = tx_pin[466];
  assign mb1_FB1_BA0_IO_017_mb1_FA2_TB1_IO_015 = tx_pin[467];
  assign mb1_FB1_BA0_IO_018_mb1_FA2_TB1_IO_032 = tx_pin[468];
  assign mb1_FB1_BA0_IO_019_mb1_FA2_TB1_IO_033 = tx_pin[469];
  assign mb1_FB1_BA0_IO_020_mb1_FA2_TB1_IO_030 = tx_pin[470];
  assign mb1_FB1_BA0_IO_021_mb1_FA2_TB1_IO_031 = tx_pin[471];
  assign mb1_FB1_BA0_IO_022_mb1_FA2_TB1_IO_008 = tx_pin[472];
  assign mb1_FB1_BA0_IO_023_mb1_FA2_TB1_IO_009 = tx_pin[473];
  assign mb1_FB1_BA0_IO_024_mb1_FA2_TB1_IO_026 = tx_pin[474];
  assign mb1_FB1_BA0_IO_025_mb1_FA2_TB1_IO_027 = tx_pin[475];
  assign mb1_FB1_BA0_IO_026_mb1_FA2_TB1_IO_024 = tx_pin[476];
  assign mb1_FB1_BA0_IO_027_mb1_FA2_TB1_IO_025 = tx_pin[477];
  assign mb1_FB1_BA0_IO_028_mb1_FA2_TB1_IO_042 = tx_pin[478];
  assign mb1_FB1_BA0_IO_029_mb1_FA2_TB1_IO_043 = tx_pin[479];
  assign mb1_FB1_BA0_IO_030_mb1_FA2_TB1_IO_020 = tx_pin[480];
  assign mb1_FB1_BA0_IO_031_mb1_FA2_TB1_IO_021 = tx_pin[481];
  assign mb1_FB1_BA0_IO_032_mb1_FA2_TB1_IO_018 = tx_pin[482];
  assign mb1_FB1_BA0_IO_033_mb1_FA2_TB1_IO_019 = tx_pin[483];
  assign mb1_FB1_BA0_IO_034_mb1_FA2_TB1_IO_036 = tx_pin[484];
  assign mb1_FB1_BA0_IO_035_mb1_FA2_TB1_IO_037 = tx_pin[485];
  assign mb1_FB1_BA0_IO_036_mb1_FA2_TB1_IO_034 = tx_pin[486];
  assign mb1_FB1_BA0_IO_037_mb1_FA2_TB1_IO_035 = tx_pin[487];
  assign mb1_FB1_BA0_IO_038_mb1_FA2_TB1_IO_052 = tx_pin[488];
  assign mb1_FB1_BA0_IO_039_mb1_FA2_TB1_IO_053 = tx_pin[489];
  assign mb1_FB1_BA0_IO_040_mb1_FA2_TB1_IO_050 = tx_pin[490];
  assign mb1_FB1_BA0_IO_041_mb1_FA2_TB1_IO_051 = tx_pin[491];
  assign mb1_FB1_BA0_IO_042_mb1_FA2_TB1_IO_028 = tx_pin[492];
  assign mb1_FB1_BA0_IO_043_mb1_FA2_TB1_IO_029 = tx_pin[493];
  assign mb1_FB1_BA0_IO_044_mb1_FA2_TB1_IO_046 = tx_pin[494];
  assign mb1_FB1_BA0_IO_045_mb1_FA2_TB1_IO_047 = tx_pin[495];
  assign mb1_FB1_BA0_IO_046_mb1_FA2_TB1_IO_044 = tx_pin[496];
  assign mb1_FB1_BA0_IO_047_mb1_FA2_TB1_IO_045 = tx_pin[497];
  assign mb1_FB1_BA0_IO_048_mb1_FA2_TB1_IO_062 = tx_pin[498];
  assign mb1_FB1_BA0_IO_049_mb1_FA2_TB1_IO_063 = tx_pin[499];
  assign mb1_FB1_BA0_IO_050_mb1_FA2_TB1_IO_040 = tx_pin[500];
  assign mb1_FB1_BA0_IO_051_mb1_FA2_TB1_IO_041 = tx_pin[501];
  assign mb1_FB1_BA0_IO_052_mb1_FA2_TB1_IO_038 = tx_pin[502];
  assign mb1_FB1_BA0_IO_053_mb1_FA2_TB1_IO_039 = tx_pin[503];
  assign mb1_FB1_BA0_IO_054_mb1_FA2_TB1_IO_056 = tx_pin[504];
  assign mb1_FB1_BA0_IO_055_mb1_FA2_TB1_IO_057 = tx_pin[505];
  assign mb1_FB1_BA0_IO_056_mb1_FA2_TB1_IO_054 = tx_pin[506];
  assign mb1_FB1_BA0_IO_057_mb1_FA2_TB1_IO_055 = tx_pin[507];
  assign mb1_FB1_BA0_IO_058_mb1_FA2_TB1_IO_072 = tx_pin[508];
  assign mb1_FB1_BA0_IO_059_mb1_FA2_TB1_IO_073 = tx_pin[509];
  assign mb1_FB1_BA0_IO_060_mb1_FA2_TB1_IO_070 = tx_pin[510];
  assign mb1_FB1_BA0_IO_061_mb1_FA2_TB1_IO_071 = tx_pin[511];
  assign mb1_FB1_BA0_IO_062_mb1_FA2_TB1_IO_048 = tx_pin[512];
  assign mb1_FB1_BA0_IO_063_mb1_FA2_TB1_IO_049 = tx_pin[513];
  assign mb1_FB1_BA0_IO_064_mb1_FA2_TB1_IO_066 = tx_pin[514];
  assign mb1_FB1_BA0_IO_065_mb1_FA2_TB1_IO_067 = tx_pin[515];
  assign mb1_FB1_BA0_IO_066_mb1_FA2_TB1_IO_064 = tx_pin[516];
  assign mb1_FB1_BA0_IO_067_mb1_FA2_TB1_IO_065 = tx_pin[517];
  assign mb1_FB1_BA0_IO_068_mb1_FA2_TB1_IO_082 = tx_pin[518];
  assign mb1_FB1_BA0_IO_069_mb1_FA2_TB1_IO_083 = tx_pin[519];
  assign mb1_FB1_BA0_IO_070_mb1_FA2_TB1_IO_060 = tx_pin[520];
  assign mb1_FB1_BA0_IO_071_mb1_FA2_TB1_IO_061 = tx_pin[521];
  assign mb1_FB1_BA0_IO_072_mb1_FA2_TB1_IO_058 = tx_pin[522];
  assign mb1_FB1_BA0_IO_073_mb1_FA2_TB1_IO_059 = tx_pin[523];
  assign mb1_FB1_BA0_IO_074_mb1_FA2_TB1_IO_076 = tx_pin[524];
  assign mb1_FB1_BA0_IO_075_mb1_FA2_TB1_IO_077 = tx_pin[525];
  assign mb1_FB1_BA0_IO_076_mb1_FA2_TB1_IO_074 = tx_pin[526];
  assign mb1_FB1_BA0_IO_077_mb1_FA2_TB1_IO_075 = tx_pin[527];
  assign mb1_FB1_BA0_IO_078_mb1_FA2_TB1_IO_092 = tx_pin[528];
  assign mb1_FB1_BA0_IO_079_mb1_FA2_TB1_IO_093 = tx_pin[529];
  assign mb1_FB1_BA0_IO_080_mb1_FA2_TB1_IO_090 = tx_pin[530];
  assign mb1_FB1_BA0_IO_081_mb1_FA2_TB1_IO_091 = tx_pin[531];
  assign mb1_FB1_BA0_IO_082_mb1_FA2_TB1_IO_068 = tx_pin[532];
  assign mb1_FB1_BA0_IO_083_mb1_FA2_TB1_IO_069 = tx_pin[533];
  assign mb1_FB1_BA0_IO_084_mb1_FA2_TB1_IO_086 = tx_pin[534];
  assign mb1_FB1_BA0_IO_085_mb1_FA2_TB1_IO_087 = tx_pin[535];
  assign mb1_FB1_BA0_IO_086_mb1_FA2_TB1_IO_084 = tx_pin[536];
  assign mb1_FB1_BA0_IO_087_mb1_FA2_TB1_IO_085 = tx_pin[537];
  assign mb1_FB1_BA0_IO_088_mb1_FA2_TB1_IO_102 = tx_pin[538];
  assign mb1_FB1_BA0_IO_089_mb1_FA2_TB1_IO_103 = tx_pin[539];
  assign mb1_FB1_BA0_IO_090_mb1_FA2_TB1_IO_080 = tx_pin[540];
  assign mb1_FB1_BA0_IO_091_mb1_FA2_TB1_IO_081 = tx_pin[541];
  assign mb1_FB1_BA0_IO_092_mb1_FA2_TB1_IO_078 = tx_pin[542];
  assign mb1_FB1_BA0_IO_093_mb1_FA2_TB1_IO_079 = tx_pin[543];
  assign mb1_FB1_BA0_IO_094_mb1_FA2_TB1_IO_096 = tx_pin[544];
  assign mb1_FB1_BA0_IO_095_mb1_FA2_TB1_IO_097 = tx_pin[545];
  assign mb1_FB1_BA0_IO_096_mb1_FA2_TB1_IO_094 = tx_pin[546];
  assign mb1_FB1_BA0_IO_097_mb1_FA2_TB1_IO_095 = tx_pin[547];
  assign mb1_FB1_BA0_IO_098_mb1_FA2_TB1_IO_112 = tx_pin[548];
  assign mb1_FB1_BA0_IO_099_mb1_FA2_TB1_IO_113 = tx_pin[549];
  assign mb1_FB1_BA0_IO_100_mb1_FA2_TB1_IO_110 = tx_pin[550];
  assign mb1_FB1_BA0_IO_101_mb1_FA2_TB1_IO_111 = tx_pin[551];
  assign mb1_FB1_BA0_IO_102_mb1_FA2_TB1_IO_088 = tx_pin[552];
  assign mb1_FB1_BA0_IO_103_mb1_FA2_TB1_IO_089 = tx_pin[553];
  assign mb1_FB1_BA0_IO_104_mb1_FA2_TB1_IO_106 = tx_pin[554];
  assign mb1_FB1_BA0_IO_105_mb1_FA2_TB1_IO_107 = tx_pin[555];
  assign mb1_FB1_BA0_IO_106_mb1_FA2_TB1_IO_104 = tx_pin[556];
  assign mb1_FB1_BA0_IO_107_mb1_FA2_TB1_IO_105 = tx_pin[557];
  assign mb1_FB1_BA0_IO_108_mb1_FA2_TB1_IO_122 = tx_pin[558];
  assign mb1_FB1_BA0_IO_109_mb1_FA2_TB1_IO_123 = tx_pin[559];
  assign mb1_FB1_BA0_IO_110_mb1_FA2_TB1_IO_100 = tx_pin[560];
  assign mb1_FB1_BA0_IO_111_mb1_FA2_TB1_IO_101 = tx_pin[561];
  assign mb1_FB1_BA0_IO_112_mb1_FA2_TB1_IO_098 = tx_pin[562];
  assign mb1_FB1_BA0_IO_113_mb1_FA2_TB1_IO_099 = tx_pin[563];
  assign mb1_FB1_BA0_IO_114_mb1_FA2_TB1_IO_116 = tx_pin[564];
  assign mb1_FB1_BA0_IO_115_mb1_FA2_TB1_IO_117 = tx_pin[565];
  assign mb1_FB1_BA0_IO_116_mb1_FA2_TB1_IO_114 = tx_pin[566];
  assign mb1_FB1_BA0_IO_117_mb1_FA2_TB1_IO_115 = tx_pin[567];
  assign mb1_FB1_BA0_IO_118_mb1_FA2_TB1_IO_132 = tx_pin[568];
  assign mb1_FB1_BA0_IO_119_mb1_FA2_TB1_IO_133 = tx_pin[569];
  assign mb1_FB1_BA0_IO_120_mb1_FA2_TB1_IO_130 = tx_pin[570];
  assign mb1_FB1_BA0_IO_121_mb1_FA2_TB1_IO_131 = tx_pin[571];
  assign mb1_FB1_BA0_IO_122_mb1_FA2_TB1_IO_108 = tx_pin[572];
  assign mb1_FB1_BA0_IO_123_mb1_FA2_TB1_IO_109 = tx_pin[573];
  assign mb1_FB1_BA0_IO_124_mb1_FA2_TB1_IO_126 = tx_pin[574];
  assign mb1_FB1_BA0_IO_125_mb1_FA2_TB1_IO_127 = tx_pin[575];
  assign mb1_FB1_BA0_IO_126_mb1_FA2_TB1_IO_124 = tx_pin[576];
  assign mb1_FB1_BA0_IO_127_mb1_FA2_TB1_IO_125 = tx_pin[577];
  assign mb1_FB1_BA0_IO_130_mb1_FA2_TB1_IO_120 = tx_pin[578];
  assign mb1_FB1_BA0_IO_131_mb1_FA2_TB1_IO_121 = tx_pin[579];
  assign mb1_FB1_BA0_IO_132_mb1_FA2_TB1_IO_118 = tx_pin[580];
  assign mb1_FB1_BA0_IO_133_mb1_FA2_TB1_IO_119 = tx_pin[581];
  assign mb1_FB1_BA0_IO_134_mb1_FA2_TB1_IO_136 = tx_pin[582];
  assign mb1_FB1_BA0_IO_136_mb1_FA2_TB1_IO_134 = tx_pin[583];
  assign mb1_FB1_BA1_CLKIO_N_0_mb1_FA2_TB0_CLKIO_N_7 = tx_pin[584];
  assign mb1_FB1_BA1_CLKIO_N_1_mb1_FA2_TB0_CLKIO_N_6 = tx_pin[585];
  assign mb1_FB1_BA1_CLKIO_N_2_mb1_FA2_TB0_CLKIO_N_4 = tx_pin[586];
  assign mb1_FB1_BA1_CLKIO_N_3_mb1_FA2_TB0_CLKIO_N_3 = tx_pin[587];
  assign mb1_FB1_BA1_CLKIO_N_4_mb1_FA2_TB0_CLKIO_N_2 = tx_pin[588];
  assign mb1_FB1_BA1_CLKIO_N_5_mb1_FA2_TB0_IO_010 = tx_pin[589];
  assign mb1_FB1_BA1_CLKIO_N_6_mb1_FA2_TB0_CLKIO_N_1 = tx_pin[590];
  assign mb1_FB1_BA1_CLKIO_N_7_mb1_FA2_TB0_CLKIO_N_0 = tx_pin[591];
  assign mb1_FB1_BA1_CLKIO_P_0_mb1_FA2_TB0_CLKIO_P_7 = tx_pin[592];
  assign mb1_FB1_BA1_CLKIO_P_1_mb1_FA2_TB0_CLKIO_P_6 = tx_pin[593];
  assign mb1_FB1_BA1_CLKIO_P_2_mb1_FA2_TB0_CLKIO_P_4 = tx_pin[594];
  assign mb1_FB1_BA1_CLKIO_P_3_mb1_FA2_TB0_CLKIO_P_3 = tx_pin[595];
  assign mb1_FB1_BA1_CLKIO_P_4_mb1_FA2_TB0_CLKIO_P_2 = tx_pin[596];
  assign mb1_FB1_BA1_CLKIO_P_5_mb1_FA2_TB0_IO_011 = tx_pin[597];
  assign mb1_FB1_BA1_CLKIO_P_6_mb1_FA2_TB0_CLKIO_P_1 = tx_pin[598];
  assign mb1_FB1_BA1_CLKIO_P_7_mb1_FA2_TB0_CLKIO_P_0 = tx_pin[599];
  assign mb1_FB1_BA1_IO_004_mb1_FA2_TB0_IO_006 = tx_pin[600];
  assign mb1_FB1_BA1_IO_005_mb1_FA2_TB0_IO_007 = tx_pin[601];
  assign mb1_FB1_BA1_IO_006_mb1_FA2_TB0_IO_004 = tx_pin[602];
  assign mb1_FB1_BA1_IO_007_mb1_FA2_TB0_IO_005 = tx_pin[603];
  assign mb1_FB1_BA1_IO_008_mb1_FA2_TB0_IO_022 = tx_pin[604];
  assign mb1_FB1_BA1_IO_009_mb1_FA2_TB0_IO_023 = tx_pin[605];
  assign mb1_FB1_BA1_IO_010_mb1_FA2_TB0_CLKIO_N_5 = tx_pin[606];
  assign mb1_FB1_BA1_IO_011_mb1_FA2_TB0_CLKIO_P_5 = tx_pin[607];
  assign mb1_FB1_BA1_IO_012_mb1_FA2_TB0_IO_012 = tx_pin[608];
  assign mb1_FB1_BA1_IO_013_mb1_FA2_TB0_IO_013 = tx_pin[609];
  assign mb1_FB1_BA1_IO_014_mb1_FA2_TB0_IO_016 = tx_pin[610];
  assign mb1_FB1_BA1_IO_015_mb1_FA2_TB0_IO_017 = tx_pin[611];
  assign mb1_FB1_BA1_IO_016_mb1_FA2_TB0_IO_014 = tx_pin[612];
  assign mb1_FB1_BA1_IO_017_mb1_FA2_TB0_IO_015 = tx_pin[613];
  assign mb1_FB1_BA1_IO_018_mb1_FA2_TB0_IO_032 = tx_pin[614];
  assign mb1_FB1_BA1_IO_019_mb1_FA2_TB0_IO_033 = tx_pin[615];
  assign mb1_FB1_BA1_IO_020_mb1_FA2_TB0_IO_030 = tx_pin[616];
  assign mb1_FB1_BA1_IO_021_mb1_FA2_TB0_IO_031 = tx_pin[617];
  assign mb1_FB1_BA1_IO_022_mb1_FA2_TB0_IO_008 = tx_pin[618];
  assign mb1_FB1_BA1_IO_023_mb1_FA2_TB0_IO_009 = tx_pin[619];
  assign mb1_FB1_BA1_IO_024_mb1_FA2_TB0_IO_026 = tx_pin[620];
  assign mb1_FB1_BA1_IO_025_mb1_FA2_TB0_IO_027 = tx_pin[621];
  assign mb1_FB1_BA1_IO_026_mb1_FA2_TB0_IO_024 = tx_pin[622];
  assign mb1_FB1_BA1_IO_027_mb1_FA2_TB0_IO_025 = tx_pin[623];
  assign mb1_FB1_BA1_IO_028_mb1_FA2_TB0_IO_042 = tx_pin[624];
  assign mb1_FB1_BA1_IO_029_mb1_FA2_TB0_IO_043 = tx_pin[625];
  assign mb1_FB1_BA1_IO_030_mb1_FA2_TB0_IO_020 = tx_pin[626];
  assign mb1_FB1_BA1_IO_031_mb1_FA2_TB0_IO_021 = tx_pin[627];
  assign mb1_FB1_BA1_IO_032_mb1_FA2_TB0_IO_018 = tx_pin[628];
  assign mb1_FB1_BA1_IO_033_mb1_FA2_TB0_IO_019 = tx_pin[629];
  assign mb1_FB1_BA1_IO_034_mb1_FA2_TB0_IO_036 = tx_pin[630];
  assign mb1_FB1_BA1_IO_035_mb1_FA2_TB0_IO_037 = tx_pin[631];
  assign mb1_FB1_BA1_IO_036_mb1_FA2_TB0_IO_034 = tx_pin[632];
  assign mb1_FB1_BA1_IO_037_mb1_FA2_TB0_IO_035 = tx_pin[633];
  assign mb1_FB1_BA1_IO_038_mb1_FA2_TB0_IO_052 = tx_pin[634];
  assign mb1_FB1_BA1_IO_039_mb1_FA2_TB0_IO_053 = tx_pin[635];
  assign mb1_FB1_BA1_IO_040_mb1_FA2_TB0_IO_050 = tx_pin[636];
  assign mb1_FB1_BA1_IO_041_mb1_FA2_TB0_IO_051 = tx_pin[637];
  assign mb1_FB1_BA1_IO_042_mb1_FA2_TB0_IO_028 = tx_pin[638];
  assign mb1_FB1_BA1_IO_043_mb1_FA2_TB0_IO_029 = tx_pin[639];
  assign mb1_FB1_BA1_IO_044_mb1_FA2_TB0_IO_046 = tx_pin[640];
  assign mb1_FB1_BA1_IO_045_mb1_FA2_TB0_IO_047 = tx_pin[641];
  assign mb1_FB1_BA1_IO_046_mb1_FA2_TB0_IO_044 = tx_pin[642];
  assign mb1_FB1_BA1_IO_047_mb1_FA2_TB0_IO_045 = tx_pin[643];
  assign mb1_FB1_BA1_IO_048_mb1_FA2_TB0_IO_062 = tx_pin[644];
  assign mb1_FB1_BA1_IO_049_mb1_FA2_TB0_IO_063 = tx_pin[645];
  assign mb1_FB1_BA1_IO_050_mb1_FA2_TB0_IO_040 = tx_pin[646];
  assign mb1_FB1_BA1_IO_051_mb1_FA2_TB0_IO_041 = tx_pin[647];
  assign mb1_FB1_BA1_IO_052_mb1_FA2_TB0_IO_038 = tx_pin[648];
  assign mb1_FB1_BA1_IO_053_mb1_FA2_TB0_IO_039 = tx_pin[649];
  assign mb1_FB1_BA1_IO_054_mb1_FA2_TB0_IO_056 = tx_pin[650];
  assign mb1_FB1_BA1_IO_055_mb1_FA2_TB0_IO_057 = tx_pin[651];
  assign mb1_FB1_BA1_IO_056_mb1_FA2_TB0_IO_054 = tx_pin[652];
  assign mb1_FB1_BA1_IO_057_mb1_FA2_TB0_IO_055 = tx_pin[653];
  assign mb1_FB1_BA1_IO_058_mb1_FA2_TB0_IO_072 = tx_pin[654];
  assign mb1_FB1_BA1_IO_059_mb1_FA2_TB0_IO_073 = tx_pin[655];
  assign mb1_FB1_BA1_IO_060_mb1_FA2_TB0_IO_070 = tx_pin[656];
  assign mb1_FB1_BA1_IO_061_mb1_FA2_TB0_IO_071 = tx_pin[657];
  assign mb1_FB1_BA1_IO_062_mb1_FA2_TB0_IO_048 = tx_pin[658];
  assign mb1_FB1_BA1_IO_063_mb1_FA2_TB0_IO_049 = tx_pin[659];
  assign mb1_FB1_BA1_IO_064_mb1_FA2_TB0_IO_066 = tx_pin[660];
  assign mb1_FB1_BA1_IO_065_mb1_FA2_TB0_IO_067 = tx_pin[661];
  assign mb1_FB1_BA1_IO_066_mb1_FA2_TB0_IO_064 = tx_pin[662];
  assign mb1_FB1_BA1_IO_067_mb1_FA2_TB0_IO_065 = tx_pin[663];
  assign mb1_FB1_BA1_IO_068_mb1_FA2_TB0_IO_082 = tx_pin[664];
  assign mb1_FB1_BA1_IO_069_mb1_FA2_TB0_IO_083 = tx_pin[665];
  assign mb1_FB1_BA1_IO_070_mb1_FA2_TB0_IO_060 = tx_pin[666];
  assign mb1_FB1_BA1_IO_071_mb1_FA2_TB0_IO_061 = tx_pin[667];
  assign mb1_FB1_BA1_IO_072_mb1_FA2_TB0_IO_058 = tx_pin[668];
  assign mb1_FB1_BA1_IO_073_mb1_FA2_TB0_IO_059 = tx_pin[669];
  assign mb1_FB1_BA1_IO_074_mb1_FA2_TB0_IO_076 = tx_pin[670];
  assign mb1_FB1_BA1_IO_075_mb1_FA2_TB0_IO_077 = tx_pin[671];
  assign mb1_FB1_BA1_IO_076_mb1_FA2_TB0_IO_074 = tx_pin[672];
  assign mb1_FB1_BA1_IO_077_mb1_FA2_TB0_IO_075 = tx_pin[673];
  assign mb1_FB1_BA1_IO_078_mb1_FA2_TB0_IO_092 = tx_pin[674];
  assign mb1_FB1_BA1_IO_079_mb1_FA2_TB0_IO_093 = tx_pin[675];
  assign mb1_FB1_BA1_IO_080_mb1_FA2_TB0_IO_090 = tx_pin[676];
  assign mb1_FB1_BA1_IO_081_mb1_FA2_TB0_IO_091 = tx_pin[677];
  assign mb1_FB1_BA1_IO_082_mb1_FA2_TB0_IO_068 = tx_pin[678];
  assign mb1_FB1_BA1_IO_083_mb1_FA2_TB0_IO_069 = tx_pin[679];
  assign mb1_FB1_BA1_IO_084_mb1_FA2_TB0_IO_086 = tx_pin[680];
  assign mb1_FB1_BA1_IO_085_mb1_FA2_TB0_IO_087 = tx_pin[681];
  assign mb1_FB1_BA1_IO_086_mb1_FA2_TB0_IO_084 = tx_pin[682];
  assign mb1_FB1_BA1_IO_087_mb1_FA2_TB0_IO_085 = tx_pin[683];
  assign mb1_FB1_BA1_IO_088_mb1_FA2_TB0_IO_102 = tx_pin[684];
  assign mb1_FB1_BA1_IO_089_mb1_FA2_TB0_IO_103 = tx_pin[685];
  assign mb1_FB1_BA1_IO_090_mb1_FA2_TB0_IO_080 = tx_pin[686];
  assign mb1_FB1_BA1_IO_091_mb1_FA2_TB0_IO_081 = tx_pin[687];
  assign mb1_FB1_BA1_IO_092_mb1_FA2_TB0_IO_078 = tx_pin[688];
  assign mb1_FB1_BA1_IO_093_mb1_FA2_TB0_IO_079 = tx_pin[689];
  assign mb1_FB1_BA1_IO_094_mb1_FA2_TB0_IO_096 = tx_pin[690];
  assign mb1_FB1_BA1_IO_095_mb1_FA2_TB0_IO_097 = tx_pin[691];
  assign mb1_FB1_BA1_IO_096_mb1_FA2_TB0_IO_094 = tx_pin[692];
  assign mb1_FB1_BA1_IO_097_mb1_FA2_TB0_IO_095 = tx_pin[693];
  assign mb1_FB1_BA1_IO_098_mb1_FA2_TB0_IO_112 = tx_pin[694];
  assign mb1_FB1_BA1_IO_099_mb1_FA2_TB0_IO_113 = tx_pin[695];
  assign mb1_FB1_BA1_IO_100_mb1_FA2_TB0_IO_110 = tx_pin[696];
  assign mb1_FB1_BA1_IO_101_mb1_FA2_TB0_IO_111 = tx_pin[697];
  assign mb1_FB1_BA1_IO_102_mb1_FA2_TB0_IO_088 = tx_pin[698];
  assign mb1_FB1_BA1_IO_103_mb1_FA2_TB0_IO_089 = tx_pin[699];
  assign mb1_FB1_BA1_IO_104_mb1_FA2_TB0_IO_106 = tx_pin[700];
  assign mb1_FB1_BA1_IO_105_mb1_FA2_TB0_IO_107 = tx_pin[701];
  assign mb1_FB1_BA1_IO_106_mb1_FA2_TB0_IO_104 = tx_pin[702];
  assign mb1_FB1_BA1_IO_107_mb1_FA2_TB0_IO_105 = tx_pin[703];
  assign mb1_FB1_BA1_IO_108_mb1_FA2_TB0_IO_122 = tx_pin[704];
  assign mb1_FB1_BA1_IO_109_mb1_FA2_TB0_IO_123 = tx_pin[705];
  assign mb1_FB1_BA1_IO_110_mb1_FA2_TB0_IO_100 = tx_pin[706];
  assign mb1_FB1_BA1_IO_111_mb1_FA2_TB0_IO_101 = tx_pin[707];
  assign mb1_FB1_BA1_IO_112_mb1_FA2_TB0_IO_098 = tx_pin[708];
  assign mb1_FB1_BA1_IO_113_mb1_FA2_TB0_IO_099 = tx_pin[709];
  assign mb1_FB1_BA1_IO_114_mb1_FA2_TB0_IO_116 = tx_pin[710];
  assign mb1_FB1_BA1_IO_115_mb1_FA2_TB0_IO_117 = tx_pin[711];
  assign mb1_FB1_BA1_IO_116_mb1_FA2_TB0_IO_114 = tx_pin[712];
  assign mb1_FB1_BA1_IO_117_mb1_FA2_TB0_IO_115 = tx_pin[713];
  assign mb1_FB1_BA1_IO_118_mb1_FA2_TB0_IO_132 = tx_pin[714];
  assign mb1_FB1_BA1_IO_119_mb1_FA2_TB0_IO_133 = tx_pin[715];
  assign mb1_FB1_BA1_IO_120_mb1_FA2_TB0_IO_130 = tx_pin[716];
  assign mb1_FB1_BA1_IO_121_mb1_FA2_TB0_IO_131 = tx_pin[717];
  assign mb1_FB1_BA1_IO_122_mb1_FA2_TB0_IO_108 = tx_pin[718];
  assign mb1_FB1_BA1_IO_123_mb1_FA2_TB0_IO_109 = tx_pin[719];
  assign mb1_FB1_BA1_IO_124_mb1_FA2_TB0_IO_126 = tx_pin[720];
  assign mb1_FB1_BA1_IO_125_mb1_FA2_TB0_IO_127 = tx_pin[721];
  assign mb1_FB1_BA1_IO_126_mb1_FA2_TB0_IO_124 = tx_pin[722];
  assign mb1_FB1_BA1_IO_127_mb1_FA2_TB0_IO_125 = tx_pin[723];
  assign mb1_FB1_BA1_IO_130_mb1_FA2_TB0_IO_120 = tx_pin[724];
  assign mb1_FB1_BA1_IO_131_mb1_FA2_TB0_IO_121 = tx_pin[725];
  assign mb1_FB1_BA1_IO_132_mb1_FA2_TB0_IO_118 = tx_pin[726];
  assign mb1_FB1_BA1_IO_133_mb1_FA2_TB0_IO_119 = tx_pin[727];
  assign mb1_FB1_BA1_IO_134_mb1_FA2_TB0_IO_136 = tx_pin[728];
  assign mb1_FB1_BA1_IO_136_mb1_FA2_TB0_IO_134 = tx_pin[729];
  assign rx_pin[292] = mb1_FA1_BA0_CLKIO_N_0_mb1_FB1_BA2_CLKIO_N_7;
  assign rx_pin[293] = mb1_FA1_BA0_CLKIO_N_1_mb1_FB1_BA2_CLKIO_N_6;
  assign rx_pin[294] = mb1_FA1_BA0_CLKIO_N_2_mb1_FB1_BA2_CLKIO_N_4;
  assign rx_pin[295] = mb1_FA1_BA0_CLKIO_N_3_mb1_FB1_BA2_CLKIO_N_3;
  assign rx_pin[296] = mb1_FA1_BA0_CLKIO_N_4_mb1_FB1_BA2_CLKIO_N_2;
  assign rx_pin[297] = mb1_FA1_BA0_CLKIO_N_5_mb1_FB1_BA2_IO_010;
  assign rx_pin[298] = mb1_FA1_BA0_CLKIO_N_6_mb1_FB1_BA2_CLKIO_N_1;
  assign rx_pin[299] = mb1_FA1_BA0_CLKIO_N_7_mb1_FB1_BA2_CLKIO_N_0;
  assign rx_pin[300] = mb1_FA1_BA0_CLKIO_P_0_mb1_FB1_BA2_CLKIO_P_7;
  assign rx_pin[301] = mb1_FA1_BA0_CLKIO_P_1_mb1_FB1_BA2_CLKIO_P_6;
  assign rx_pin[302] = mb1_FA1_BA0_CLKIO_P_2_mb1_FB1_BA2_CLKIO_P_4;
  assign rx_pin[303] = mb1_FA1_BA0_CLKIO_P_3_mb1_FB1_BA2_CLKIO_P_3;
  assign rx_pin[304] = mb1_FA1_BA0_CLKIO_P_4_mb1_FB1_BA2_CLKIO_P_2;
  assign rx_pin[305] = mb1_FA1_BA0_CLKIO_P_5_mb1_FB1_BA2_IO_011;
  assign rx_pin[306] = mb1_FA1_BA0_CLKIO_P_6_mb1_FB1_BA2_CLKIO_P_1;
  assign rx_pin[307] = mb1_FA1_BA0_CLKIO_P_7_mb1_FB1_BA2_CLKIO_P_0;
  assign rx_pin[308] = mb1_FA1_BA0_IO_004_mb1_FB1_BA2_IO_006;
  assign rx_pin[309] = mb1_FA1_BA0_IO_005_mb1_FB1_BA2_IO_007;
  assign rx_pin[310] = mb1_FA1_BA0_IO_006_mb1_FB1_BA2_IO_004;
  assign rx_pin[311] = mb1_FA1_BA0_IO_007_mb1_FB1_BA2_IO_005;
  assign rx_pin[312] = mb1_FA1_BA0_IO_008_mb1_FB1_BA2_IO_022;
  assign rx_pin[313] = mb1_FA1_BA0_IO_009_mb1_FB1_BA2_IO_023;
  assign rx_pin[314] = mb1_FA1_BA0_IO_010_mb1_FB1_BA2_CLKIO_N_5;
  assign rx_pin[315] = mb1_FA1_BA0_IO_011_mb1_FB1_BA2_CLKIO_P_5;
  assign rx_pin[316] = mb1_FA1_BA0_IO_012_mb1_FB1_BA2_IO_012;
  assign rx_pin[317] = mb1_FA1_BA0_IO_013_mb1_FB1_BA2_IO_013;
  assign rx_pin[318] = mb1_FA1_BA0_IO_014_mb1_FB1_BA2_IO_016;
  assign rx_pin[319] = mb1_FA1_BA0_IO_015_mb1_FB1_BA2_IO_017;
  assign rx_pin[320] = mb1_FA1_BA0_IO_016_mb1_FB1_BA2_IO_014;
  assign rx_pin[321] = mb1_FA1_BA0_IO_017_mb1_FB1_BA2_IO_015;
  assign rx_pin[322] = mb1_FA1_BA0_IO_018_mb1_FB1_BA2_IO_032;
  assign rx_pin[323] = mb1_FA1_BA0_IO_019_mb1_FB1_BA2_IO_033;
  assign rx_pin[324] = mb1_FA1_BA0_IO_020_mb1_FB1_BA2_IO_030;
  assign rx_pin[325] = mb1_FA1_BA0_IO_021_mb1_FB1_BA2_IO_031;
  assign rx_pin[326] = mb1_FA1_BA0_IO_022_mb1_FB1_BA2_IO_008;
  assign rx_pin[327] = mb1_FA1_BA0_IO_023_mb1_FB1_BA2_IO_009;
  assign rx_pin[328] = mb1_FA1_BA0_IO_024_mb1_FB1_BA2_IO_026;
  assign rx_pin[329] = mb1_FA1_BA0_IO_025_mb1_FB1_BA2_IO_027;
  assign rx_pin[330] = mb1_FA1_BA0_IO_026_mb1_FB1_BA2_IO_024;
  assign rx_pin[331] = mb1_FA1_BA0_IO_027_mb1_FB1_BA2_IO_025;
  assign rx_pin[332] = mb1_FA1_BA0_IO_028_mb1_FB1_BA2_IO_042;
  assign rx_pin[333] = mb1_FA1_BA0_IO_029_mb1_FB1_BA2_IO_043;
  assign rx_pin[334] = mb1_FA1_BA0_IO_030_mb1_FB1_BA2_IO_020;
  assign rx_pin[335] = mb1_FA1_BA0_IO_031_mb1_FB1_BA2_IO_021;
  assign rx_pin[336] = mb1_FA1_BA0_IO_032_mb1_FB1_BA2_IO_018;
  assign rx_pin[337] = mb1_FA1_BA0_IO_033_mb1_FB1_BA2_IO_019;
  assign rx_pin[338] = mb1_FA1_BA0_IO_034_mb1_FB1_BA2_IO_036;
  assign rx_pin[339] = mb1_FA1_BA0_IO_035_mb1_FB1_BA2_IO_037;
  assign rx_pin[340] = mb1_FA1_BA0_IO_036_mb1_FB1_BA2_IO_034;
  assign rx_pin[341] = mb1_FA1_BA0_IO_037_mb1_FB1_BA2_IO_035;
  assign rx_pin[342] = mb1_FA1_BA0_IO_038_mb1_FB1_BA2_IO_052;
  assign rx_pin[343] = mb1_FA1_BA0_IO_039_mb1_FB1_BA2_IO_053;
  assign rx_pin[344] = mb1_FA1_BA0_IO_040_mb1_FB1_BA2_IO_050;
  assign rx_pin[345] = mb1_FA1_BA0_IO_041_mb1_FB1_BA2_IO_051;
  assign rx_pin[346] = mb1_FA1_BA0_IO_042_mb1_FB1_BA2_IO_028;
  assign rx_pin[347] = mb1_FA1_BA0_IO_043_mb1_FB1_BA2_IO_029;
  assign rx_pin[348] = mb1_FA1_BA0_IO_044_mb1_FB1_BA2_IO_046;
  assign rx_pin[349] = mb1_FA1_BA0_IO_045_mb1_FB1_BA2_IO_047;
  assign rx_pin[350] = mb1_FA1_BA0_IO_046_mb1_FB1_BA2_IO_044;
  assign rx_pin[351] = mb1_FA1_BA0_IO_047_mb1_FB1_BA2_IO_045;
  assign rx_pin[352] = mb1_FA1_BA0_IO_048_mb1_FB1_BA2_IO_062;
  assign rx_pin[353] = mb1_FA1_BA0_IO_049_mb1_FB1_BA2_IO_063;
  assign rx_pin[354] = mb1_FA1_BA0_IO_050_mb1_FB1_BA2_IO_040;
  assign rx_pin[355] = mb1_FA1_BA0_IO_051_mb1_FB1_BA2_IO_041;
  assign rx_pin[356] = mb1_FA1_BA0_IO_052_mb1_FB1_BA2_IO_038;
  assign rx_pin[357] = mb1_FA1_BA0_IO_053_mb1_FB1_BA2_IO_039;
  assign rx_pin[358] = mb1_FA1_BA0_IO_054_mb1_FB1_BA2_IO_056;
  assign rx_pin[359] = mb1_FA1_BA0_IO_055_mb1_FB1_BA2_IO_057;
  assign rx_pin[360] = mb1_FA1_BA0_IO_056_mb1_FB1_BA2_IO_054;
  assign rx_pin[361] = mb1_FA1_BA0_IO_057_mb1_FB1_BA2_IO_055;
  assign rx_pin[362] = mb1_FA1_BA0_IO_058_mb1_FB1_BA2_IO_072;
  assign rx_pin[363] = mb1_FA1_BA0_IO_059_mb1_FB1_BA2_IO_073;
  assign rx_pin[364] = mb1_FA1_BA0_IO_060_mb1_FB1_BA2_IO_070;
  assign rx_pin[365] = mb1_FA1_BA0_IO_061_mb1_FB1_BA2_IO_071;
  assign rx_pin[366] = mb1_FA1_BA0_IO_062_mb1_FB1_BA2_IO_048;
  assign rx_pin[367] = mb1_FA1_BA0_IO_063_mb1_FB1_BA2_IO_049;
  assign rx_pin[368] = mb1_FA1_BA0_IO_064_mb1_FB1_BA2_IO_066;
  assign rx_pin[369] = mb1_FA1_BA0_IO_065_mb1_FB1_BA2_IO_067;
  assign rx_pin[370] = mb1_FA1_BA0_IO_066_mb1_FB1_BA2_IO_064;
  assign rx_pin[371] = mb1_FA1_BA0_IO_067_mb1_FB1_BA2_IO_065;
  assign rx_pin[372] = mb1_FA1_BA0_IO_068_mb1_FB1_BA2_IO_082;
  assign rx_pin[373] = mb1_FA1_BA0_IO_069_mb1_FB1_BA2_IO_083;
  assign rx_pin[374] = mb1_FA1_BA0_IO_070_mb1_FB1_BA2_IO_060;
  assign rx_pin[375] = mb1_FA1_BA0_IO_071_mb1_FB1_BA2_IO_061;
  assign rx_pin[376] = mb1_FA1_BA0_IO_072_mb1_FB1_BA2_IO_058;
  assign rx_pin[377] = mb1_FA1_BA0_IO_073_mb1_FB1_BA2_IO_059;
  assign rx_pin[378] = mb1_FA1_BA0_IO_074_mb1_FB1_BA2_IO_076;
  assign rx_pin[379] = mb1_FA1_BA0_IO_075_mb1_FB1_BA2_IO_077;
  assign rx_pin[380] = mb1_FA1_BA0_IO_076_mb1_FB1_BA2_IO_074;
  assign rx_pin[381] = mb1_FA1_BA0_IO_077_mb1_FB1_BA2_IO_075;
  assign rx_pin[382] = mb1_FA1_BA0_IO_078_mb1_FB1_BA2_IO_092;
  assign rx_pin[383] = mb1_FA1_BA0_IO_079_mb1_FB1_BA2_IO_093;
  assign rx_pin[384] = mb1_FA1_BA0_IO_080_mb1_FB1_BA2_IO_090;
  assign rx_pin[385] = mb1_FA1_BA0_IO_081_mb1_FB1_BA2_IO_091;
  assign rx_pin[386] = mb1_FA1_BA0_IO_082_mb1_FB1_BA2_IO_068;
  assign rx_pin[387] = mb1_FA1_BA0_IO_083_mb1_FB1_BA2_IO_069;
  assign rx_pin[388] = mb1_FA1_BA0_IO_084_mb1_FB1_BA2_IO_086;
  assign rx_pin[389] = mb1_FA1_BA0_IO_085_mb1_FB1_BA2_IO_087;
  assign rx_pin[390] = mb1_FA1_BA0_IO_086_mb1_FB1_BA2_IO_084;
  assign rx_pin[391] = mb1_FA1_BA0_IO_087_mb1_FB1_BA2_IO_085;
  assign rx_pin[392] = mb1_FA1_BA0_IO_088_mb1_FB1_BA2_IO_102;
  assign rx_pin[393] = mb1_FA1_BA0_IO_089_mb1_FB1_BA2_IO_103;
  assign rx_pin[394] = mb1_FA1_BA0_IO_090_mb1_FB1_BA2_IO_080;
  assign rx_pin[395] = mb1_FA1_BA0_IO_091_mb1_FB1_BA2_IO_081;
  assign rx_pin[396] = mb1_FA1_BA0_IO_092_mb1_FB1_BA2_IO_078;
  assign rx_pin[397] = mb1_FA1_BA0_IO_093_mb1_FB1_BA2_IO_079;
  assign rx_pin[398] = mb1_FA1_BA0_IO_094_mb1_FB1_BA2_IO_096;
  assign rx_pin[399] = mb1_FA1_BA0_IO_095_mb1_FB1_BA2_IO_097;
  assign rx_pin[400] = mb1_FA1_BA0_IO_096_mb1_FB1_BA2_IO_094;
  assign rx_pin[401] = mb1_FA1_BA0_IO_097_mb1_FB1_BA2_IO_095;
  assign rx_pin[402] = mb1_FA1_BA0_IO_098_mb1_FB1_BA2_IO_112;
  assign rx_pin[403] = mb1_FA1_BA0_IO_099_mb1_FB1_BA2_IO_113;
  assign rx_pin[404] = mb1_FA1_BA0_IO_100_mb1_FB1_BA2_IO_110;
  assign rx_pin[405] = mb1_FA1_BA0_IO_101_mb1_FB1_BA2_IO_111;
  assign rx_pin[406] = mb1_FA1_BA0_IO_102_mb1_FB1_BA2_IO_088;
  assign rx_pin[407] = mb1_FA1_BA0_IO_103_mb1_FB1_BA2_IO_089;
  assign rx_pin[408] = mb1_FA1_BA0_IO_104_mb1_FB1_BA2_IO_106;
  assign rx_pin[409] = mb1_FA1_BA0_IO_105_mb1_FB1_BA2_IO_107;
  assign rx_pin[410] = mb1_FA1_BA0_IO_106_mb1_FB1_BA2_IO_104;
  assign rx_pin[411] = mb1_FA1_BA0_IO_107_mb1_FB1_BA2_IO_105;
  assign rx_pin[412] = mb1_FA1_BA0_IO_108_mb1_FB1_BA2_IO_122;
  assign rx_pin[413] = mb1_FA1_BA0_IO_109_mb1_FB1_BA2_IO_123;
  assign rx_pin[414] = mb1_FA1_BA0_IO_110_mb1_FB1_BA2_IO_100;
  assign rx_pin[415] = mb1_FA1_BA0_IO_111_mb1_FB1_BA2_IO_101;
  assign rx_pin[416] = mb1_FA1_BA0_IO_112_mb1_FB1_BA2_IO_098;
  assign rx_pin[417] = mb1_FA1_BA0_IO_113_mb1_FB1_BA2_IO_099;
  assign rx_pin[418] = mb1_FA1_BA0_IO_114_mb1_FB1_BA2_IO_116;
  assign rx_pin[419] = mb1_FA1_BA0_IO_115_mb1_FB1_BA2_IO_117;
  assign rx_pin[420] = mb1_FA1_BA0_IO_116_mb1_FB1_BA2_IO_114;
  assign rx_pin[421] = mb1_FA1_BA0_IO_117_mb1_FB1_BA2_IO_115;
  assign rx_pin[422] = mb1_FA1_BA0_IO_118_mb1_FB1_BA2_IO_132;
  assign rx_pin[423] = mb1_FA1_BA0_IO_119_mb1_FB1_BA2_IO_133;
  assign rx_pin[424] = mb1_FA1_BA0_IO_120_mb1_FB1_BA2_IO_130;
  assign rx_pin[425] = mb1_FA1_BA0_IO_121_mb1_FB1_BA2_IO_131;
  assign rx_pin[426] = mb1_FA1_BA0_IO_122_mb1_FB1_BA2_IO_108;
  assign rx_pin[427] = mb1_FA1_BA0_IO_123_mb1_FB1_BA2_IO_109;
  assign rx_pin[428] = mb1_FA1_BA0_IO_124_mb1_FB1_BA2_IO_126;
  assign rx_pin[429] = mb1_FA1_BA0_IO_125_mb1_FB1_BA2_IO_127;
  assign rx_pin[430] = mb1_FA1_BA0_IO_126_mb1_FB1_BA2_IO_124;
  assign rx_pin[431] = mb1_FA1_BA0_IO_127_mb1_FB1_BA2_IO_125;
  assign rx_pin[432] = mb1_FA1_BA0_IO_130_mb1_FB1_BA2_IO_120;
  assign rx_pin[433] = mb1_FA1_BA0_IO_131_mb1_FB1_BA2_IO_121;
  assign rx_pin[434] = mb1_FA1_BA0_IO_132_mb1_FB1_BA2_IO_118;
  assign rx_pin[435] = mb1_FA1_BA0_IO_133_mb1_FB1_BA2_IO_119;
  assign rx_pin[436] = mb1_FA1_BA0_IO_134_mb1_FB1_BA2_IO_136;
  assign rx_pin[437] = mb1_FA1_BA0_IO_136_mb1_FB1_BA2_IO_134;
  assign rx_pin[438] = mb1_FA1_BA2_CLKIO_N_0_mb1_FB1_BB0_CLKIO_N_7;
  assign rx_pin[439] = mb1_FA1_BA2_CLKIO_N_1_mb1_FB1_BB0_CLKIO_N_6;
  assign rx_pin[440] = mb1_FA1_BA2_CLKIO_N_2_mb1_FB1_BB0_CLKIO_N_4;
  assign rx_pin[441] = mb1_FA1_BA2_CLKIO_N_3_mb1_FB1_BB0_CLKIO_N_3;
  assign rx_pin[442] = mb1_FA1_BA2_CLKIO_N_4_mb1_FB1_BB0_CLKIO_N_2;
  assign rx_pin[443] = mb1_FA1_BA2_CLKIO_N_5_mb1_FB1_BB0_IO_010;
  assign rx_pin[444] = mb1_FA1_BA2_CLKIO_N_6_mb1_FB1_BB0_CLKIO_N_1;
  assign rx_pin[445] = mb1_FA1_BA2_CLKIO_N_7_mb1_FB1_BB0_CLKIO_N_0;
  assign rx_pin[446] = mb1_FA1_BA2_CLKIO_P_0_mb1_FB1_BB0_CLKIO_P_7;
  assign rx_pin[447] = mb1_FA1_BA2_CLKIO_P_1_mb1_FB1_BB0_CLKIO_P_6;
  assign rx_pin[448] = mb1_FA1_BA2_CLKIO_P_2_mb1_FB1_BB0_CLKIO_P_4;
  assign rx_pin[449] = mb1_FA1_BA2_CLKIO_P_3_mb1_FB1_BB0_CLKIO_P_3;
  assign rx_pin[450] = mb1_FA1_BA2_CLKIO_P_4_mb1_FB1_BB0_CLKIO_P_2;
  assign rx_pin[451] = mb1_FA1_BA2_CLKIO_P_5_mb1_FB1_BB0_IO_011;
  assign rx_pin[452] = mb1_FA1_BA2_CLKIO_P_6_mb1_FB1_BB0_CLKIO_P_1;
  assign rx_pin[453] = mb1_FA1_BA2_CLKIO_P_7_mb1_FB1_BB0_CLKIO_P_0;
  assign rx_pin[454] = mb1_FA1_BA2_IO_004_mb1_FB1_BB0_IO_006;
  assign rx_pin[455] = mb1_FA1_BA2_IO_005_mb1_FB1_BB0_IO_007;
  assign rx_pin[456] = mb1_FA1_BA2_IO_006_mb1_FB1_BB0_IO_004;
  assign rx_pin[457] = mb1_FA1_BA2_IO_007_mb1_FB1_BB0_IO_005;
  assign rx_pin[458] = mb1_FA1_BA2_IO_008_mb1_FB1_BB0_IO_022;
  assign rx_pin[459] = mb1_FA1_BA2_IO_009_mb1_FB1_BB0_IO_023;
  assign rx_pin[460] = mb1_FA1_BA2_IO_010_mb1_FB1_BB0_CLKIO_N_5;
  assign rx_pin[461] = mb1_FA1_BA2_IO_011_mb1_FB1_BB0_CLKIO_P_5;
  assign rx_pin[462] = mb1_FA1_BA2_IO_012_mb1_FB1_BB0_IO_012;
  assign rx_pin[463] = mb1_FA1_BA2_IO_013_mb1_FB1_BB0_IO_013;
  assign rx_pin[464] = mb1_FA1_BA2_IO_014_mb1_FB1_BB0_IO_016;
  assign rx_pin[465] = mb1_FA1_BA2_IO_015_mb1_FB1_BB0_IO_017;
  assign rx_pin[466] = mb1_FA1_BA2_IO_016_mb1_FB1_BB0_IO_014;
  assign rx_pin[467] = mb1_FA1_BA2_IO_017_mb1_FB1_BB0_IO_015;
  assign rx_pin[468] = mb1_FA1_BA2_IO_018_mb1_FB1_BB0_IO_032;
  assign rx_pin[469] = mb1_FA1_BA2_IO_019_mb1_FB1_BB0_IO_033;
  assign rx_pin[470] = mb1_FA1_BA2_IO_020_mb1_FB1_BB0_IO_030;
  assign rx_pin[471] = mb1_FA1_BA2_IO_021_mb1_FB1_BB0_IO_031;
  assign rx_pin[472] = mb1_FA1_BA2_IO_022_mb1_FB1_BB0_IO_008;
  assign rx_pin[473] = mb1_FA1_BA2_IO_023_mb1_FB1_BB0_IO_009;
  assign rx_pin[474] = mb1_FA1_BA2_IO_024_mb1_FB1_BB0_IO_026;
  assign rx_pin[475] = mb1_FA1_BA2_IO_025_mb1_FB1_BB0_IO_027;
  assign rx_pin[476] = mb1_FA1_BA2_IO_026_mb1_FB1_BB0_IO_024;
  assign rx_pin[477] = mb1_FA1_BA2_IO_027_mb1_FB1_BB0_IO_025;
  assign rx_pin[478] = mb1_FA1_BA2_IO_028_mb1_FB1_BB0_IO_042;
  assign rx_pin[479] = mb1_FA1_BA2_IO_029_mb1_FB1_BB0_IO_043;
  assign rx_pin[480] = mb1_FA1_BA2_IO_030_mb1_FB1_BB0_IO_020;
  assign rx_pin[481] = mb1_FA1_BA2_IO_031_mb1_FB1_BB0_IO_021;
  assign rx_pin[482] = mb1_FA1_BA2_IO_032_mb1_FB1_BB0_IO_018;
  assign rx_pin[483] = mb1_FA1_BA2_IO_033_mb1_FB1_BB0_IO_019;
  assign rx_pin[484] = mb1_FA1_BA2_IO_034_mb1_FB1_BB0_IO_036;
  assign rx_pin[485] = mb1_FA1_BA2_IO_035_mb1_FB1_BB0_IO_037;
  assign rx_pin[486] = mb1_FA1_BA2_IO_036_mb1_FB1_BB0_IO_034;
  assign rx_pin[487] = mb1_FA1_BA2_IO_037_mb1_FB1_BB0_IO_035;
  assign rx_pin[488] = mb1_FA1_BA2_IO_038_mb1_FB1_BB0_IO_052;
  assign rx_pin[489] = mb1_FA1_BA2_IO_039_mb1_FB1_BB0_IO_053;
  assign rx_pin[490] = mb1_FA1_BA2_IO_040_mb1_FB1_BB0_IO_050;
  assign rx_pin[491] = mb1_FA1_BA2_IO_041_mb1_FB1_BB0_IO_051;
  assign rx_pin[492] = mb1_FA1_BA2_IO_042_mb1_FB1_BB0_IO_028;
  assign rx_pin[493] = mb1_FA1_BA2_IO_043_mb1_FB1_BB0_IO_029;
  assign rx_pin[494] = mb1_FA1_BA2_IO_044_mb1_FB1_BB0_IO_046;
  assign rx_pin[495] = mb1_FA1_BA2_IO_045_mb1_FB1_BB0_IO_047;
  assign rx_pin[496] = mb1_FA1_BA2_IO_046_mb1_FB1_BB0_IO_044;
  assign rx_pin[497] = mb1_FA1_BA2_IO_047_mb1_FB1_BB0_IO_045;
  assign rx_pin[498] = mb1_FA1_BA2_IO_048_mb1_FB1_BB0_IO_062;
  assign rx_pin[499] = mb1_FA1_BA2_IO_049_mb1_FB1_BB0_IO_063;
  assign rx_pin[500] = mb1_FA1_BA2_IO_050_mb1_FB1_BB0_IO_040;
  assign rx_pin[501] = mb1_FA1_BA2_IO_051_mb1_FB1_BB0_IO_041;
  assign rx_pin[502] = mb1_FA1_BA2_IO_052_mb1_FB1_BB0_IO_038;
  assign rx_pin[503] = mb1_FA1_BA2_IO_053_mb1_FB1_BB0_IO_039;
  assign rx_pin[504] = mb1_FA1_BA2_IO_054_mb1_FB1_BB0_IO_056;
  assign rx_pin[505] = mb1_FA1_BA2_IO_055_mb1_FB1_BB0_IO_057;
  assign rx_pin[506] = mb1_FA1_BA2_IO_056_mb1_FB1_BB0_IO_054;
  assign rx_pin[507] = mb1_FA1_BA2_IO_057_mb1_FB1_BB0_IO_055;
  assign rx_pin[508] = mb1_FA1_BA2_IO_058_mb1_FB1_BB0_IO_072;
  assign rx_pin[509] = mb1_FA1_BA2_IO_059_mb1_FB1_BB0_IO_073;
  assign rx_pin[510] = mb1_FA1_BA2_IO_060_mb1_FB1_BB0_IO_070;
  assign rx_pin[511] = mb1_FA1_BA2_IO_061_mb1_FB1_BB0_IO_071;
  assign rx_pin[512] = mb1_FA1_BA2_IO_062_mb1_FB1_BB0_IO_048;
  assign rx_pin[513] = mb1_FA1_BA2_IO_063_mb1_FB1_BB0_IO_049;
  assign rx_pin[514] = mb1_FA1_BA2_IO_064_mb1_FB1_BB0_IO_066;
  assign rx_pin[515] = mb1_FA1_BA2_IO_065_mb1_FB1_BB0_IO_067;
  assign rx_pin[516] = mb1_FA1_BA2_IO_066_mb1_FB1_BB0_IO_064;
  assign rx_pin[517] = mb1_FA1_BA2_IO_067_mb1_FB1_BB0_IO_065;
  assign rx_pin[518] = mb1_FA1_BA2_IO_068_mb1_FB1_BB0_IO_082;
  assign rx_pin[519] = mb1_FA1_BA2_IO_069_mb1_FB1_BB0_IO_083;
  assign rx_pin[520] = mb1_FA1_BA2_IO_070_mb1_FB1_BB0_IO_060;
  assign rx_pin[521] = mb1_FA1_BA2_IO_071_mb1_FB1_BB0_IO_061;
  assign rx_pin[522] = mb1_FA1_BA2_IO_072_mb1_FB1_BB0_IO_058;
  assign rx_pin[523] = mb1_FA1_BA2_IO_073_mb1_FB1_BB0_IO_059;
  assign rx_pin[524] = mb1_FA1_BA2_IO_074_mb1_FB1_BB0_IO_076;
  assign rx_pin[525] = mb1_FA1_BA2_IO_075_mb1_FB1_BB0_IO_077;
  assign rx_pin[526] = mb1_FA1_BA2_IO_076_mb1_FB1_BB0_IO_074;
  assign rx_pin[527] = mb1_FA1_BA2_IO_077_mb1_FB1_BB0_IO_075;
  assign rx_pin[528] = mb1_FA1_BA2_IO_078_mb1_FB1_BB0_IO_092;
  assign rx_pin[529] = mb1_FA1_BA2_IO_079_mb1_FB1_BB0_IO_093;
  assign rx_pin[530] = mb1_FA1_BA2_IO_080_mb1_FB1_BB0_IO_090;
  assign rx_pin[531] = mb1_FA1_BA2_IO_081_mb1_FB1_BB0_IO_091;
  assign rx_pin[532] = mb1_FA1_BA2_IO_082_mb1_FB1_BB0_IO_068;
  assign rx_pin[533] = mb1_FA1_BA2_IO_083_mb1_FB1_BB0_IO_069;
  assign rx_pin[534] = mb1_FA1_BA2_IO_084_mb1_FB1_BB0_IO_086;
  assign rx_pin[535] = mb1_FA1_BA2_IO_085_mb1_FB1_BB0_IO_087;
  assign rx_pin[536] = mb1_FA1_BA2_IO_086_mb1_FB1_BB0_IO_084;
  assign rx_pin[537] = mb1_FA1_BA2_IO_087_mb1_FB1_BB0_IO_085;
  assign rx_pin[538] = mb1_FA1_BA2_IO_088_mb1_FB1_BB0_IO_102;
  assign rx_pin[539] = mb1_FA1_BA2_IO_089_mb1_FB1_BB0_IO_103;
  assign rx_pin[540] = mb1_FA1_BA2_IO_090_mb1_FB1_BB0_IO_080;
  assign rx_pin[541] = mb1_FA1_BA2_IO_091_mb1_FB1_BB0_IO_081;
  assign rx_pin[542] = mb1_FA1_BA2_IO_092_mb1_FB1_BB0_IO_078;
  assign rx_pin[543] = mb1_FA1_BA2_IO_093_mb1_FB1_BB0_IO_079;
  assign rx_pin[544] = mb1_FA1_BA2_IO_094_mb1_FB1_BB0_IO_096;
  assign rx_pin[545] = mb1_FA1_BA2_IO_095_mb1_FB1_BB0_IO_097;
  assign rx_pin[546] = mb1_FA1_BA2_IO_096_mb1_FB1_BB0_IO_094;
  assign rx_pin[547] = mb1_FA1_BA2_IO_097_mb1_FB1_BB0_IO_095;
  assign rx_pin[548] = mb1_FA1_BA2_IO_098_mb1_FB1_BB0_IO_112;
  assign rx_pin[549] = mb1_FA1_BA2_IO_099_mb1_FB1_BB0_IO_113;
  assign rx_pin[550] = mb1_FA1_BA2_IO_100_mb1_FB1_BB0_IO_110;
  assign rx_pin[551] = mb1_FA1_BA2_IO_101_mb1_FB1_BB0_IO_111;
  assign rx_pin[552] = mb1_FA1_BA2_IO_102_mb1_FB1_BB0_IO_088;
  assign rx_pin[553] = mb1_FA1_BA2_IO_103_mb1_FB1_BB0_IO_089;
  assign rx_pin[554] = mb1_FA1_BA2_IO_104_mb1_FB1_BB0_IO_106;
  assign rx_pin[555] = mb1_FA1_BA2_IO_105_mb1_FB1_BB0_IO_107;
  assign rx_pin[556] = mb1_FA1_BA2_IO_106_mb1_FB1_BB0_IO_104;
  assign rx_pin[557] = mb1_FA1_BA2_IO_107_mb1_FB1_BB0_IO_105;
  assign rx_pin[558] = mb1_FA1_BA2_IO_108_mb1_FB1_BB0_IO_122;
  assign rx_pin[559] = mb1_FA1_BA2_IO_109_mb1_FB1_BB0_IO_123;
  assign rx_pin[560] = mb1_FA1_BA2_IO_110_mb1_FB1_BB0_IO_100;
  assign rx_pin[561] = mb1_FA1_BA2_IO_111_mb1_FB1_BB0_IO_101;
  assign rx_pin[562] = mb1_FA1_BA2_IO_112_mb1_FB1_BB0_IO_098;
  assign rx_pin[563] = mb1_FA1_BA2_IO_113_mb1_FB1_BB0_IO_099;
  assign rx_pin[564] = mb1_FA1_BA2_IO_114_mb1_FB1_BB0_IO_116;
  assign rx_pin[565] = mb1_FA1_BA2_IO_115_mb1_FB1_BB0_IO_117;
  assign rx_pin[566] = mb1_FA1_BA2_IO_116_mb1_FB1_BB0_IO_114;
  assign rx_pin[567] = mb1_FA1_BA2_IO_117_mb1_FB1_BB0_IO_115;
  assign rx_pin[568] = mb1_FA1_BA2_IO_118_mb1_FB1_BB0_IO_132;
  assign rx_pin[569] = mb1_FA1_BA2_IO_119_mb1_FB1_BB0_IO_133;
  assign rx_pin[570] = mb1_FA1_BA2_IO_120_mb1_FB1_BB0_IO_130;
  assign rx_pin[571] = mb1_FA1_BA2_IO_121_mb1_FB1_BB0_IO_131;
  assign rx_pin[572] = mb1_FA1_BA2_IO_122_mb1_FB1_BB0_IO_108;
  assign rx_pin[573] = mb1_FA1_BA2_IO_123_mb1_FB1_BB0_IO_109;
  assign rx_pin[574] = mb1_FA1_BA2_IO_124_mb1_FB1_BB0_IO_126;
  assign rx_pin[575] = mb1_FA1_BA2_IO_125_mb1_FB1_BB0_IO_127;
  assign rx_pin[576] = mb1_FA1_BA2_IO_126_mb1_FB1_BB0_IO_124;
  assign rx_pin[577] = mb1_FA1_BA2_IO_127_mb1_FB1_BB0_IO_125;
  assign rx_pin[578] = mb1_FA1_BA2_IO_130_mb1_FB1_BB0_IO_120;
  assign rx_pin[579] = mb1_FA1_BA2_IO_131_mb1_FB1_BB0_IO_121;
  assign rx_pin[580] = mb1_FA1_BA2_IO_132_mb1_FB1_BB0_IO_118;
  assign rx_pin[581] = mb1_FA1_BA2_IO_133_mb1_FB1_BB0_IO_119;
  assign rx_pin[582] = mb1_FA1_BA2_IO_134_mb1_FB1_BB0_IO_136;
  assign rx_pin[583] = mb1_FA1_BA2_IO_136_mb1_FB1_BB0_IO_134;
  assign rx_pin[584] = mb1_FA1_TB1_CLKIO_N_0_mb1_FB1_BB1_CLKIO_N_7;
  assign rx_pin[585] = mb1_FA1_TB1_CLKIO_N_1_mb1_FB1_BB1_CLKIO_N_6;
  assign rx_pin[586] = mb1_FA1_TB1_CLKIO_N_2_mb1_FB1_BB1_CLKIO_N_4;
  assign rx_pin[587] = mb1_FA1_TB1_CLKIO_N_3_mb1_FB1_BB1_CLKIO_N_3;
  assign rx_pin[588] = mb1_FA1_TB1_CLKIO_N_4_mb1_FB1_BB1_CLKIO_N_2;
  assign rx_pin[589] = mb1_FA1_TB1_CLKIO_N_5_mb1_FB1_BB1_IO_010;
  assign rx_pin[590] = mb1_FA1_TB1_CLKIO_N_6_mb1_FB1_BB1_CLKIO_N_1;
  assign rx_pin[591] = mb1_FA1_TB1_CLKIO_N_7_mb1_FB1_BB1_CLKIO_N_0;
  assign rx_pin[592] = mb1_FA1_TB1_CLKIO_P_0_mb1_FB1_BB1_CLKIO_P_7;
  assign rx_pin[593] = mb1_FA1_TB1_CLKIO_P_1_mb1_FB1_BB1_CLKIO_P_6;
  assign rx_pin[594] = mb1_FA1_TB1_CLKIO_P_2_mb1_FB1_BB1_CLKIO_P_4;
  assign rx_pin[595] = mb1_FA1_TB1_CLKIO_P_3_mb1_FB1_BB1_CLKIO_P_3;
  assign rx_pin[596] = mb1_FA1_TB1_CLKIO_P_4_mb1_FB1_BB1_CLKIO_P_2;
  assign rx_pin[597] = mb1_FA1_TB1_CLKIO_P_5_mb1_FB1_BB1_IO_011;
  assign rx_pin[598] = mb1_FA1_TB1_CLKIO_P_6_mb1_FB1_BB1_CLKIO_P_1;
  assign rx_pin[599] = mb1_FA1_TB1_CLKIO_P_7_mb1_FB1_BB1_CLKIO_P_0;
  assign rx_pin[600] = mb1_FA1_TB1_IO_004_mb1_FB1_BB1_IO_006;
  assign rx_pin[601] = mb1_FA1_TB1_IO_005_mb1_FB1_BB1_IO_007;
  assign rx_pin[602] = mb1_FA1_TB1_IO_006_mb1_FB1_BB1_IO_004;
  assign rx_pin[603] = mb1_FA1_TB1_IO_007_mb1_FB1_BB1_IO_005;
  assign rx_pin[604] = mb1_FA1_TB1_IO_008_mb1_FB1_BB1_IO_022;
  assign rx_pin[605] = mb1_FA1_TB1_IO_009_mb1_FB1_BB1_IO_023;
  assign rx_pin[606] = mb1_FA1_TB1_IO_010_mb1_FB1_BB1_CLKIO_N_5;
  assign rx_pin[607] = mb1_FA1_TB1_IO_011_mb1_FB1_BB1_CLKIO_P_5;
  assign rx_pin[608] = mb1_FA1_TB1_IO_012_mb1_FB1_BB1_IO_012;
  assign rx_pin[609] = mb1_FA1_TB1_IO_013_mb1_FB1_BB1_IO_013;
  assign rx_pin[610] = mb1_FA1_TB1_IO_014_mb1_FB1_BB1_IO_016;
  assign rx_pin[611] = mb1_FA1_TB1_IO_015_mb1_FB1_BB1_IO_017;
  assign rx_pin[612] = mb1_FA1_TB1_IO_016_mb1_FB1_BB1_IO_014;
  assign rx_pin[613] = mb1_FA1_TB1_IO_017_mb1_FB1_BB1_IO_015;
  assign rx_pin[614] = mb1_FA1_TB1_IO_018_mb1_FB1_BB1_IO_032;
  assign rx_pin[615] = mb1_FA1_TB1_IO_019_mb1_FB1_BB1_IO_033;
  assign rx_pin[616] = mb1_FA1_TB1_IO_020_mb1_FB1_BB1_IO_030;
  assign rx_pin[617] = mb1_FA1_TB1_IO_021_mb1_FB1_BB1_IO_031;
  assign rx_pin[618] = mb1_FA1_TB1_IO_022_mb1_FB1_BB1_IO_008;
  assign rx_pin[619] = mb1_FA1_TB1_IO_023_mb1_FB1_BB1_IO_009;
  assign rx_pin[620] = mb1_FA1_TB1_IO_024_mb1_FB1_BB1_IO_026;
  assign rx_pin[621] = mb1_FA1_TB1_IO_025_mb1_FB1_BB1_IO_027;
  assign rx_pin[622] = mb1_FA1_TB1_IO_026_mb1_FB1_BB1_IO_024;
  assign rx_pin[623] = mb1_FA1_TB1_IO_027_mb1_FB1_BB1_IO_025;
  assign rx_pin[624] = mb1_FA1_TB1_IO_028_mb1_FB1_BB1_IO_042;
  assign rx_pin[625] = mb1_FA1_TB1_IO_029_mb1_FB1_BB1_IO_043;
  assign rx_pin[626] = mb1_FA1_TB1_IO_030_mb1_FB1_BB1_IO_020;
  assign rx_pin[627] = mb1_FA1_TB1_IO_031_mb1_FB1_BB1_IO_021;
  assign rx_pin[628] = mb1_FA1_TB1_IO_032_mb1_FB1_BB1_IO_018;
  assign rx_pin[629] = mb1_FA1_TB1_IO_033_mb1_FB1_BB1_IO_019;
  assign rx_pin[630] = mb1_FA1_TB1_IO_034_mb1_FB1_BB1_IO_036;
  assign rx_pin[631] = mb1_FA1_TB1_IO_035_mb1_FB1_BB1_IO_037;
  assign rx_pin[632] = mb1_FA1_TB1_IO_036_mb1_FB1_BB1_IO_034;
  assign rx_pin[633] = mb1_FA1_TB1_IO_037_mb1_FB1_BB1_IO_035;
  assign rx_pin[634] = mb1_FA1_TB1_IO_038_mb1_FB1_BB1_IO_052;
  assign rx_pin[635] = mb1_FA1_TB1_IO_039_mb1_FB1_BB1_IO_053;
  assign rx_pin[636] = mb1_FA1_TB1_IO_040_mb1_FB1_BB1_IO_050;
  assign rx_pin[637] = mb1_FA1_TB1_IO_041_mb1_FB1_BB1_IO_051;
  assign rx_pin[638] = mb1_FA1_TB1_IO_042_mb1_FB1_BB1_IO_028;
  assign rx_pin[639] = mb1_FA1_TB1_IO_043_mb1_FB1_BB1_IO_029;
  assign rx_pin[640] = mb1_FA1_TB1_IO_044_mb1_FB1_BB1_IO_046;
  assign rx_pin[641] = mb1_FA1_TB1_IO_045_mb1_FB1_BB1_IO_047;
  assign rx_pin[642] = mb1_FA1_TB1_IO_046_mb1_FB1_BB1_IO_044;
  assign rx_pin[643] = mb1_FA1_TB1_IO_047_mb1_FB1_BB1_IO_045;
  assign rx_pin[644] = mb1_FA1_TB1_IO_048_mb1_FB1_BB1_IO_062;
  assign rx_pin[645] = mb1_FA1_TB1_IO_049_mb1_FB1_BB1_IO_063;
  assign rx_pin[646] = mb1_FA1_TB1_IO_050_mb1_FB1_BB1_IO_040;
  assign rx_pin[647] = mb1_FA1_TB1_IO_051_mb1_FB1_BB1_IO_041;
  assign rx_pin[648] = mb1_FA1_TB1_IO_052_mb1_FB1_BB1_IO_038;
  assign rx_pin[649] = mb1_FA1_TB1_IO_053_mb1_FB1_BB1_IO_039;
  assign rx_pin[650] = mb1_FA1_TB1_IO_054_mb1_FB1_BB1_IO_056;
  assign rx_pin[651] = mb1_FA1_TB1_IO_055_mb1_FB1_BB1_IO_057;
  assign rx_pin[652] = mb1_FA1_TB1_IO_056_mb1_FB1_BB1_IO_054;
  assign rx_pin[653] = mb1_FA1_TB1_IO_057_mb1_FB1_BB1_IO_055;
  assign rx_pin[654] = mb1_FA1_TB1_IO_058_mb1_FB1_BB1_IO_072;
  assign rx_pin[655] = mb1_FA1_TB1_IO_059_mb1_FB1_BB1_IO_073;
  assign rx_pin[656] = mb1_FA1_TB1_IO_060_mb1_FB1_BB1_IO_070;
  assign rx_pin[657] = mb1_FA1_TB1_IO_061_mb1_FB1_BB1_IO_071;
  assign rx_pin[658] = mb1_FA1_TB1_IO_062_mb1_FB1_BB1_IO_048;
  assign rx_pin[659] = mb1_FA1_TB1_IO_063_mb1_FB1_BB1_IO_049;
  assign rx_pin[660] = mb1_FA1_TB1_IO_064_mb1_FB1_BB1_IO_066;
  assign rx_pin[661] = mb1_FA1_TB1_IO_065_mb1_FB1_BB1_IO_067;
  assign rx_pin[662] = mb1_FA1_TB1_IO_066_mb1_FB1_BB1_IO_064;
  assign rx_pin[663] = mb1_FA1_TB1_IO_067_mb1_FB1_BB1_IO_065;
  assign rx_pin[664] = mb1_FA1_TB1_IO_068_mb1_FB1_BB1_IO_082;
  assign rx_pin[665] = mb1_FA1_TB1_IO_069_mb1_FB1_BB1_IO_083;
  assign rx_pin[666] = mb1_FA1_TB1_IO_070_mb1_FB1_BB1_IO_060;
  assign rx_pin[667] = mb1_FA1_TB1_IO_071_mb1_FB1_BB1_IO_061;
  assign rx_pin[668] = mb1_FA1_TB1_IO_072_mb1_FB1_BB1_IO_058;
  assign rx_pin[669] = mb1_FA1_TB1_IO_073_mb1_FB1_BB1_IO_059;
  assign rx_pin[670] = mb1_FA1_TB1_IO_074_mb1_FB1_BB1_IO_076;
  assign rx_pin[671] = mb1_FA1_TB1_IO_075_mb1_FB1_BB1_IO_077;
  assign rx_pin[672] = mb1_FA1_TB1_IO_076_mb1_FB1_BB1_IO_074;
  assign rx_pin[673] = mb1_FA1_TB1_IO_077_mb1_FB1_BB1_IO_075;
  assign rx_pin[674] = mb1_FA1_TB1_IO_078_mb1_FB1_BB1_IO_092;
  assign rx_pin[675] = mb1_FA1_TB1_IO_079_mb1_FB1_BB1_IO_093;
  assign rx_pin[676] = mb1_FA1_TB1_IO_080_mb1_FB1_BB1_IO_090;
  assign rx_pin[677] = mb1_FA1_TB1_IO_081_mb1_FB1_BB1_IO_091;
  assign rx_pin[678] = mb1_FA1_TB1_IO_082_mb1_FB1_BB1_IO_068;
  assign rx_pin[679] = mb1_FA1_TB1_IO_083_mb1_FB1_BB1_IO_069;
  assign rx_pin[680] = mb1_FA1_TB1_IO_084_mb1_FB1_BB1_IO_086;
  assign rx_pin[681] = mb1_FA1_TB1_IO_085_mb1_FB1_BB1_IO_087;
  assign rx_pin[682] = mb1_FA1_TB1_IO_086_mb1_FB1_BB1_IO_084;
  assign rx_pin[683] = mb1_FA1_TB1_IO_087_mb1_FB1_BB1_IO_085;
  assign rx_pin[684] = mb1_FA1_TB1_IO_088_mb1_FB1_BB1_IO_102;
  assign rx_pin[685] = mb1_FA1_TB1_IO_089_mb1_FB1_BB1_IO_103;
  assign rx_pin[686] = mb1_FA1_TB1_IO_090_mb1_FB1_BB1_IO_080;
  assign rx_pin[687] = mb1_FA1_TB1_IO_091_mb1_FB1_BB1_IO_081;
  assign rx_pin[688] = mb1_FA1_TB1_IO_092_mb1_FB1_BB1_IO_078;
  assign rx_pin[689] = mb1_FA1_TB1_IO_093_mb1_FB1_BB1_IO_079;
  assign rx_pin[690] = mb1_FA1_TB1_IO_094_mb1_FB1_BB1_IO_096;
  assign rx_pin[691] = mb1_FA1_TB1_IO_095_mb1_FB1_BB1_IO_097;
  assign rx_pin[692] = mb1_FA1_TB1_IO_096_mb1_FB1_BB1_IO_094;
  assign rx_pin[693] = mb1_FA1_TB1_IO_097_mb1_FB1_BB1_IO_095;
  assign rx_pin[694] = mb1_FA1_TB1_IO_098_mb1_FB1_BB1_IO_112;
  assign rx_pin[695] = mb1_FA1_TB1_IO_099_mb1_FB1_BB1_IO_113;
  assign rx_pin[696] = mb1_FA1_TB1_IO_100_mb1_FB1_BB1_IO_110;
  assign rx_pin[697] = mb1_FA1_TB1_IO_101_mb1_FB1_BB1_IO_111;
  assign rx_pin[698] = mb1_FA1_TB1_IO_102_mb1_FB1_BB1_IO_088;
  assign rx_pin[699] = mb1_FA1_TB1_IO_103_mb1_FB1_BB1_IO_089;
  assign rx_pin[700] = mb1_FA1_TB1_IO_104_mb1_FB1_BB1_IO_106;
  assign rx_pin[701] = mb1_FA1_TB1_IO_105_mb1_FB1_BB1_IO_107;
  assign rx_pin[702] = mb1_FA1_TB1_IO_106_mb1_FB1_BB1_IO_104;
  assign rx_pin[703] = mb1_FA1_TB1_IO_107_mb1_FB1_BB1_IO_105;
  assign rx_pin[704] = mb1_FA1_TB1_IO_108_mb1_FB1_BB1_IO_122;
  assign rx_pin[705] = mb1_FA1_TB1_IO_109_mb1_FB1_BB1_IO_123;
  assign rx_pin[706] = mb1_FA1_TB1_IO_110_mb1_FB1_BB1_IO_100;
  assign rx_pin[707] = mb1_FA1_TB1_IO_111_mb1_FB1_BB1_IO_101;
  assign rx_pin[708] = mb1_FA1_TB1_IO_112_mb1_FB1_BB1_IO_098;
  assign rx_pin[709] = mb1_FA1_TB1_IO_113_mb1_FB1_BB1_IO_099;
  assign rx_pin[710] = mb1_FA1_TB1_IO_114_mb1_FB1_BB1_IO_116;
  assign rx_pin[711] = mb1_FA1_TB1_IO_115_mb1_FB1_BB1_IO_117;
  assign rx_pin[712] = mb1_FA1_TB1_IO_116_mb1_FB1_BB1_IO_114;
  assign rx_pin[713] = mb1_FA1_TB1_IO_117_mb1_FB1_BB1_IO_115;
  assign rx_pin[714] = mb1_FA1_TB1_IO_118_mb1_FB1_BB1_IO_132;
  assign rx_pin[715] = mb1_FA1_TB1_IO_119_mb1_FB1_BB1_IO_133;
  assign rx_pin[716] = mb1_FA1_TB1_IO_120_mb1_FB1_BB1_IO_130;
  assign rx_pin[717] = mb1_FA1_TB1_IO_121_mb1_FB1_BB1_IO_131;
  assign rx_pin[718] = mb1_FA1_TB1_IO_122_mb1_FB1_BB1_IO_108;
  assign rx_pin[719] = mb1_FA1_TB1_IO_123_mb1_FB1_BB1_IO_109;
  assign rx_pin[720] = mb1_FA1_TB1_IO_124_mb1_FB1_BB1_IO_126;
  assign rx_pin[721] = mb1_FA1_TB1_IO_125_mb1_FB1_BB1_IO_127;
  assign rx_pin[722] = mb1_FA1_TB1_IO_126_mb1_FB1_BB1_IO_124;
  assign rx_pin[723] = mb1_FA1_TB1_IO_127_mb1_FB1_BB1_IO_125;
  assign rx_pin[724] = mb1_FA1_TB1_IO_130_mb1_FB1_BB1_IO_120;
  assign rx_pin[725] = mb1_FA1_TB1_IO_131_mb1_FB1_BB1_IO_121;
  assign rx_pin[726] = mb1_FA1_TB1_IO_132_mb1_FB1_BB1_IO_118;
  assign rx_pin[727] = mb1_FA1_TB1_IO_133_mb1_FB1_BB1_IO_119;
  assign rx_pin[728] = mb1_FA1_TB1_IO_134_mb1_FB1_BB1_IO_136;
  assign rx_pin[729] = mb1_FA1_TB1_IO_136_mb1_FB1_BB1_IO_134;
  assign rx_pin[730] = mb1_FA1_BB0_CLKIO_N_0_mb1_FB1_BB2_CLKIO_N_7;
  assign rx_pin[731] = mb1_FA1_BB0_CLKIO_N_1_mb1_FB1_BB2_CLKIO_N_6;
  assign rx_pin[732] = mb1_FA1_BB0_CLKIO_N_2_mb1_FB1_BB2_CLKIO_N_4;
  assign rx_pin[733] = mb1_FA1_BB0_CLKIO_N_3_mb1_FB1_BB2_CLKIO_N_3;
  assign rx_pin[734] = mb1_FA1_BB0_CLKIO_N_4_mb1_FB1_BB2_CLKIO_N_2;
  assign rx_pin[735] = mb1_FA1_BB0_CLKIO_N_5_mb1_FB1_BB2_IO_010;
  assign rx_pin[736] = mb1_FA1_BB0_CLKIO_N_6_mb1_FB1_BB2_CLKIO_N_1;
  assign rx_pin[737] = mb1_FA1_BB0_CLKIO_N_7_mb1_FB1_BB2_CLKIO_N_0;
  assign rx_pin[738] = mb1_FA1_BB0_CLKIO_P_0_mb1_FB1_BB2_CLKIO_P_7;
  assign rx_pin[739] = mb1_FA1_BB0_CLKIO_P_1_mb1_FB1_BB2_CLKIO_P_6;
  assign rx_pin[740] = mb1_FA1_BB0_CLKIO_P_2_mb1_FB1_BB2_CLKIO_P_4;
  assign rx_pin[741] = mb1_FA1_BB0_CLKIO_P_3_mb1_FB1_BB2_CLKIO_P_3;
  assign rx_pin[742] = mb1_FA1_BB0_CLKIO_P_4_mb1_FB1_BB2_CLKIO_P_2;
  assign rx_pin[743] = mb1_FA1_BB0_CLKIO_P_5_mb1_FB1_BB2_IO_011;
  assign rx_pin[744] = mb1_FA1_BB0_CLKIO_P_6_mb1_FB1_BB2_CLKIO_P_1;
  assign rx_pin[745] = mb1_FA1_BB0_CLKIO_P_7_mb1_FB1_BB2_CLKIO_P_0;
  assign rx_pin[746] = mb1_FA1_BB0_IO_004_mb1_FB1_BB2_IO_006;
  assign rx_pin[747] = mb1_FA1_BB0_IO_005_mb1_FB1_BB2_IO_007;
  assign rx_pin[748] = mb1_FA1_BB0_IO_006_mb1_FB1_BB2_IO_004;
  assign rx_pin[749] = mb1_FA1_BB0_IO_007_mb1_FB1_BB2_IO_005;
  assign rx_pin[750] = mb1_FA1_BB0_IO_008_mb1_FB1_BB2_IO_022;
  assign rx_pin[751] = mb1_FA1_BB0_IO_009_mb1_FB1_BB2_IO_023;
  assign rx_pin[752] = mb1_FA1_BB0_IO_010_mb1_FB1_BB2_CLKIO_N_5;
  assign rx_pin[753] = mb1_FA1_BB0_IO_011_mb1_FB1_BB2_CLKIO_P_5;
  assign rx_pin[754] = mb1_FA1_BB0_IO_012_mb1_FB1_BB2_IO_012;
  assign rx_pin[755] = mb1_FA1_BB0_IO_013_mb1_FB1_BB2_IO_013;
  assign rx_pin[756] = mb1_FA1_BB0_IO_014_mb1_FB1_BB2_IO_016;
  assign rx_pin[757] = mb1_FA1_BB0_IO_015_mb1_FB1_BB2_IO_017;
  assign rx_pin[758] = mb1_FA1_BB0_IO_016_mb1_FB1_BB2_IO_014;
  assign rx_pin[759] = mb1_FA1_BB0_IO_017_mb1_FB1_BB2_IO_015;
  assign rx_pin[760] = mb1_FA1_BB0_IO_018_mb1_FB1_BB2_IO_032;
  assign rx_pin[761] = mb1_FA1_BB0_IO_019_mb1_FB1_BB2_IO_033;
  assign rx_pin[762] = mb1_FA1_BB0_IO_020_mb1_FB1_BB2_IO_030;
  assign rx_pin[763] = mb1_FA1_BB0_IO_021_mb1_FB1_BB2_IO_031;
  assign rx_pin[764] = mb1_FA1_BB0_IO_022_mb1_FB1_BB2_IO_008;
  assign rx_pin[765] = mb1_FA1_BB0_IO_023_mb1_FB1_BB2_IO_009;
  assign rx_pin[766] = mb1_FA1_BB0_IO_024_mb1_FB1_BB2_IO_026;
  assign rx_pin[767] = mb1_FA1_BB0_IO_025_mb1_FB1_BB2_IO_027;
  assign rx_pin[768] = mb1_FA1_BB0_IO_026_mb1_FB1_BB2_IO_024;
  assign rx_pin[769] = mb1_FA1_BB0_IO_027_mb1_FB1_BB2_IO_025;
  assign rx_pin[770] = mb1_FA1_BB0_IO_028_mb1_FB1_BB2_IO_042;
  assign rx_pin[771] = mb1_FA1_BB0_IO_029_mb1_FB1_BB2_IO_043;
  assign rx_pin[772] = mb1_FA1_BB0_IO_030_mb1_FB1_BB2_IO_020;
  assign rx_pin[773] = mb1_FA1_BB0_IO_031_mb1_FB1_BB2_IO_021;
  assign rx_pin[774] = mb1_FA1_BB0_IO_032_mb1_FB1_BB2_IO_018;
  assign rx_pin[775] = mb1_FA1_BB0_IO_033_mb1_FB1_BB2_IO_019;
  assign rx_pin[776] = mb1_FA1_BB0_IO_034_mb1_FB1_BB2_IO_036;
  assign rx_pin[777] = mb1_FA1_BB0_IO_035_mb1_FB1_BB2_IO_037;
  assign rx_pin[778] = mb1_FA1_BB0_IO_036_mb1_FB1_BB2_IO_034;
  assign rx_pin[779] = mb1_FA1_BB0_IO_037_mb1_FB1_BB2_IO_035;
  assign rx_pin[780] = mb1_FA1_BB0_IO_038_mb1_FB1_BB2_IO_052;
  assign rx_pin[781] = mb1_FA1_BB0_IO_039_mb1_FB1_BB2_IO_053;
  assign rx_pin[782] = mb1_FA1_BB0_IO_040_mb1_FB1_BB2_IO_050;
  assign rx_pin[783] = mb1_FA1_BB0_IO_041_mb1_FB1_BB2_IO_051;
  assign rx_pin[784] = mb1_FA1_BB0_IO_042_mb1_FB1_BB2_IO_028;
  assign rx_pin[785] = mb1_FA1_BB0_IO_043_mb1_FB1_BB2_IO_029;
  assign rx_pin[786] = mb1_FA1_BB0_IO_044_mb1_FB1_BB2_IO_046;
  assign rx_pin[787] = mb1_FA1_BB0_IO_045_mb1_FB1_BB2_IO_047;
  assign rx_pin[788] = mb1_FA1_BB0_IO_046_mb1_FB1_BB2_IO_044;
  assign rx_pin[789] = mb1_FA1_BB0_IO_047_mb1_FB1_BB2_IO_045;
  assign rx_pin[790] = mb1_FA1_BB0_IO_048_mb1_FB1_BB2_IO_062;
  assign rx_pin[791] = mb1_FA1_BB0_IO_049_mb1_FB1_BB2_IO_063;
  assign rx_pin[792] = mb1_FA1_BB0_IO_050_mb1_FB1_BB2_IO_040;
  assign rx_pin[793] = mb1_FA1_BB0_IO_051_mb1_FB1_BB2_IO_041;
  assign rx_pin[794] = mb1_FA1_BB0_IO_052_mb1_FB1_BB2_IO_038;
  assign rx_pin[795] = mb1_FA1_BB0_IO_053_mb1_FB1_BB2_IO_039;
  assign rx_pin[796] = mb1_FA1_BB0_IO_054_mb1_FB1_BB2_IO_056;
  assign rx_pin[797] = mb1_FA1_BB0_IO_055_mb1_FB1_BB2_IO_057;
  assign rx_pin[798] = mb1_FA1_BB0_IO_056_mb1_FB1_BB2_IO_054;
  assign rx_pin[799] = mb1_FA1_BB0_IO_057_mb1_FB1_BB2_IO_055;
  assign rx_pin[800] = mb1_FA1_BB0_IO_058_mb1_FB1_BB2_IO_072;
  assign rx_pin[801] = mb1_FA1_BB0_IO_059_mb1_FB1_BB2_IO_073;
  assign rx_pin[802] = mb1_FA1_BB0_IO_060_mb1_FB1_BB2_IO_070;
  assign rx_pin[803] = mb1_FA1_BB0_IO_061_mb1_FB1_BB2_IO_071;
  assign rx_pin[804] = mb1_FA1_BB0_IO_062_mb1_FB1_BB2_IO_048;
  assign rx_pin[805] = mb1_FA1_BB0_IO_063_mb1_FB1_BB2_IO_049;
  assign rx_pin[806] = mb1_FA1_BB0_IO_064_mb1_FB1_BB2_IO_066;
  assign rx_pin[807] = mb1_FA1_BB0_IO_065_mb1_FB1_BB2_IO_067;
  assign rx_pin[808] = mb1_FA1_BB0_IO_066_mb1_FB1_BB2_IO_064;
  assign rx_pin[809] = mb1_FA1_BB0_IO_067_mb1_FB1_BB2_IO_065;
  assign rx_pin[810] = mb1_FA1_BB0_IO_068_mb1_FB1_BB2_IO_082;
  assign rx_pin[811] = mb1_FA1_BB0_IO_069_mb1_FB1_BB2_IO_083;
  assign rx_pin[812] = mb1_FA1_BB0_IO_070_mb1_FB1_BB2_IO_060;
  assign rx_pin[813] = mb1_FA1_BB0_IO_071_mb1_FB1_BB2_IO_061;
  assign rx_pin[814] = mb1_FA1_BB0_IO_072_mb1_FB1_BB2_IO_058;
  assign rx_pin[815] = mb1_FA1_BB0_IO_073_mb1_FB1_BB2_IO_059;
  assign rx_pin[816] = mb1_FA1_BB0_IO_074_mb1_FB1_BB2_IO_076;
  assign rx_pin[817] = mb1_FA1_BB0_IO_075_mb1_FB1_BB2_IO_077;
  assign rx_pin[818] = mb1_FA1_BB0_IO_076_mb1_FB1_BB2_IO_074;
  assign rx_pin[819] = mb1_FA1_BB0_IO_077_mb1_FB1_BB2_IO_075;
  assign rx_pin[820] = mb1_FA1_BB0_IO_078_mb1_FB1_BB2_IO_092;
  assign rx_pin[821] = mb1_FA1_BB0_IO_079_mb1_FB1_BB2_IO_093;
  assign rx_pin[822] = mb1_FA1_BB0_IO_080_mb1_FB1_BB2_IO_090;
  assign rx_pin[823] = mb1_FA1_BB0_IO_081_mb1_FB1_BB2_IO_091;
  assign rx_pin[824] = mb1_FA1_BB0_IO_082_mb1_FB1_BB2_IO_068;
  assign rx_pin[825] = mb1_FA1_BB0_IO_083_mb1_FB1_BB2_IO_069;
  assign rx_pin[826] = mb1_FA1_BB0_IO_084_mb1_FB1_BB2_IO_086;
  assign rx_pin[827] = mb1_FA1_BB0_IO_085_mb1_FB1_BB2_IO_087;
  assign rx_pin[828] = mb1_FA1_BB0_IO_086_mb1_FB1_BB2_IO_084;
  assign rx_pin[829] = mb1_FA1_BB0_IO_087_mb1_FB1_BB2_IO_085;
  assign rx_pin[830] = mb1_FA1_BB0_IO_088_mb1_FB1_BB2_IO_102;
  assign rx_pin[831] = mb1_FA1_BB0_IO_089_mb1_FB1_BB2_IO_103;
  assign rx_pin[832] = mb1_FA1_BB0_IO_090_mb1_FB1_BB2_IO_080;
  assign rx_pin[833] = mb1_FA1_BB0_IO_091_mb1_FB1_BB2_IO_081;
  assign rx_pin[834] = mb1_FA1_BB0_IO_092_mb1_FB1_BB2_IO_078;
  assign rx_pin[835] = mb1_FA1_BB0_IO_093_mb1_FB1_BB2_IO_079;
  assign rx_pin[836] = mb1_FA1_BB0_IO_094_mb1_FB1_BB2_IO_096;
  assign rx_pin[837] = mb1_FA1_BB0_IO_095_mb1_FB1_BB2_IO_097;
  assign rx_pin[838] = mb1_FA1_BB0_IO_096_mb1_FB1_BB2_IO_094;
  assign rx_pin[839] = mb1_FA1_BB0_IO_097_mb1_FB1_BB2_IO_095;
  assign rx_pin[840] = mb1_FA1_BB0_IO_098_mb1_FB1_BB2_IO_112;
  assign rx_pin[841] = mb1_FA1_BB0_IO_099_mb1_FB1_BB2_IO_113;
  assign rx_pin[842] = mb1_FA1_BB0_IO_100_mb1_FB1_BB2_IO_110;
  assign rx_pin[843] = mb1_FA1_BB0_IO_101_mb1_FB1_BB2_IO_111;
  assign rx_pin[844] = mb1_FA1_BB0_IO_102_mb1_FB1_BB2_IO_088;
  assign rx_pin[845] = mb1_FA1_BB0_IO_103_mb1_FB1_BB2_IO_089;
  assign rx_pin[846] = mb1_FA1_BB0_IO_104_mb1_FB1_BB2_IO_106;
  assign rx_pin[847] = mb1_FA1_BB0_IO_105_mb1_FB1_BB2_IO_107;
  assign rx_pin[848] = mb1_FA1_BB0_IO_106_mb1_FB1_BB2_IO_104;
  assign rx_pin[849] = mb1_FA1_BB0_IO_107_mb1_FB1_BB2_IO_105;
  assign rx_pin[850] = mb1_FA1_BB0_IO_108_mb1_FB1_BB2_IO_122;
  assign rx_pin[851] = mb1_FA1_BB0_IO_109_mb1_FB1_BB2_IO_123;
  assign rx_pin[852] = mb1_FA1_BB0_IO_110_mb1_FB1_BB2_IO_100;
  assign rx_pin[853] = mb1_FA1_BB0_IO_111_mb1_FB1_BB2_IO_101;
  assign rx_pin[854] = mb1_FA1_BB0_IO_112_mb1_FB1_BB2_IO_098;
  assign rx_pin[855] = mb1_FA1_BB0_IO_113_mb1_FB1_BB2_IO_099;
  assign rx_pin[856] = mb1_FA1_BB0_IO_114_mb1_FB1_BB2_IO_116;
  assign rx_pin[857] = mb1_FA1_BB0_IO_115_mb1_FB1_BB2_IO_117;
  assign rx_pin[858] = mb1_FA1_BB0_IO_116_mb1_FB1_BB2_IO_114;
  assign rx_pin[859] = mb1_FA1_BB0_IO_117_mb1_FB1_BB2_IO_115;
  assign rx_pin[860] = mb1_FA1_BB0_IO_118_mb1_FB1_BB2_IO_132;
  assign rx_pin[861] = mb1_FA1_BB0_IO_119_mb1_FB1_BB2_IO_133;
  assign rx_pin[862] = mb1_FA1_BB0_IO_120_mb1_FB1_BB2_IO_130;
  assign rx_pin[863] = mb1_FA1_BB0_IO_121_mb1_FB1_BB2_IO_131;
  assign rx_pin[864] = mb1_FA1_BB0_IO_122_mb1_FB1_BB2_IO_108;
  assign rx_pin[865] = mb1_FA1_BB0_IO_123_mb1_FB1_BB2_IO_109;
  assign rx_pin[866] = mb1_FA1_BB0_IO_124_mb1_FB1_BB2_IO_126;
  assign rx_pin[867] = mb1_FA1_BB0_IO_125_mb1_FB1_BB2_IO_127;
  assign rx_pin[868] = mb1_FA1_BB0_IO_126_mb1_FB1_BB2_IO_124;
  assign rx_pin[869] = mb1_FA1_BB0_IO_127_mb1_FB1_BB2_IO_125;
  assign rx_pin[870] = mb1_FA1_BB0_IO_130_mb1_FB1_BB2_IO_120;
  assign rx_pin[871] = mb1_FA1_BB0_IO_131_mb1_FB1_BB2_IO_121;
  assign rx_pin[872] = mb1_FA1_BB0_IO_132_mb1_FB1_BB2_IO_118;
  assign rx_pin[873] = mb1_FA1_BB0_IO_133_mb1_FB1_BB2_IO_119;
  assign rx_pin[874] = mb1_FA1_BB0_IO_134_mb1_FB1_BB2_IO_136;
  assign rx_pin[875] = mb1_FA1_BB0_IO_136_mb1_FB1_BB2_IO_134;

  dbst # (
    .DEVICE             ( "XVUP"   ),
    .TX_PINS            ( TX_PINS               ),
    .RX_PINS            ( RX_PINS               ),
    .DIFF_ENABLED       ( 0 ),
    .USE_CLK_INPUT_BUFG ( USE_CLK_INPUT_BUFG    )
  ) U_DBST (
    .tx_pin        ( tx_pin      ),
    .tx_pin_p      (             ),
    .tx_pin_n      (             ),
    .rx_pin        ( rx_pin      ),
    .rx_pin_p      ( '0          ),
    .rx_pin_n      ( '0          ),
    .clk_p         ( CLK_P[1:0]  ),
    .clk_n         ( CLK_N[1:0]  ),
    .sync_p        ( SYNC_P[1:0] ),
    .sync_n        ( SYNC_N[1:0] ),
    .dmbi_f2h_o    ( DMBI_F2H    ),
    .dmbi_h2f_i    ( DMBI_H2F    )
  );
  
endmodule
