// Unpublished work. Copyright 2022 Siemens                         
// This material contains trade secrets or otherwise                
// confidential information owned by Siemens Industry Software Inc. 
// or its affiliates (collectively, "SISW"), or its licensors.      
// Access to and use of this information is strictly limited as     
// set forth in the Customer's applicable agreements with SISW.     
// This file was generated by profpga_brdgen version 14.0 
//   on Fri Dec 15 16:10:02 2023 

`timescale 1 ps / 1 ps

// Disable implicit declaration of wires
`default_nettype none

module top_fpga_mb1fa1
   (
    input  wire [7:0]  CLK_N,
    input  wire [7:0]  CLK_P,
    input  wire [7:0]  SYNC_N,
    input  wire [7:0]  SYNC_P,
    output wire [3:0]  SRC_CLK_N,
    output wire [3:0]  SRC_CLK_P,
    output wire [3:0]  SRC_SYNC_N,
    output wire [3:0]  SRC_SYNC_P,
    output wire [19:0] DMBI_F2H,
    input  wire [19:0] DMBI_H2F,
    output wire        mb1_FA1_TA1_CLKIO_N_0_mb1_FB1_TA2_CLKIO_N_7,
    output wire        mb1_FA1_TA1_CLKIO_N_1_mb1_FB1_TA2_CLKIO_N_6,
    output wire        mb1_FA1_TA1_CLKIO_N_2_mb1_FB1_TA2_CLKIO_N_4,
    output wire        mb1_FA1_TA1_CLKIO_N_3_mb1_FB1_TA2_CLKIO_N_3,
    output wire        mb1_FA1_TA1_CLKIO_N_4_mb1_FB1_TA2_CLKIO_N_2,
    output wire        mb1_FA1_TA1_CLKIO_N_5_mb1_FB1_TA2_IO_010,
    output wire        mb1_FA1_TA1_CLKIO_N_6_mb1_FB1_TA2_CLKIO_N_1,
    output wire        mb1_FA1_TA1_CLKIO_N_7_mb1_FB1_TA2_CLKIO_N_0,
    output wire        mb1_FA1_TA1_CLKIO_P_0_mb1_FB1_TA2_CLKIO_P_7,
    output wire        mb1_FA1_TA1_CLKIO_P_1_mb1_FB1_TA2_CLKIO_P_6,
    output wire        mb1_FA1_TA1_CLKIO_P_2_mb1_FB1_TA2_CLKIO_P_4,
    output wire        mb1_FA1_TA1_CLKIO_P_3_mb1_FB1_TA2_CLKIO_P_3,
    output wire        mb1_FA1_TA1_CLKIO_P_4_mb1_FB1_TA2_CLKIO_P_2,
    output wire        mb1_FA1_TA1_CLKIO_P_5_mb1_FB1_TA2_IO_011,
    output wire        mb1_FA1_TA1_CLKIO_P_6_mb1_FB1_TA2_CLKIO_P_1,
    output wire        mb1_FA1_TA1_CLKIO_P_7_mb1_FB1_TA2_CLKIO_P_0,
    output wire        mb1_FA1_TA1_IO_004_mb1_FB1_TA2_IO_006,
    output wire        mb1_FA1_TA1_IO_005_mb1_FB1_TA2_IO_007,
    output wire        mb1_FA1_TA1_IO_006_mb1_FB1_TA2_IO_004,
    output wire        mb1_FA1_TA1_IO_007_mb1_FB1_TA2_IO_005,
    output wire        mb1_FA1_TA1_IO_008_mb1_FB1_TA2_IO_022,
    output wire        mb1_FA1_TA1_IO_009_mb1_FB1_TA2_IO_023,
    output wire        mb1_FA1_TA1_IO_010_mb1_FB1_TA2_CLKIO_N_5,
    output wire        mb1_FA1_TA1_IO_011_mb1_FB1_TA2_CLKIO_P_5,
    output wire        mb1_FA1_TA1_IO_012_mb1_FB1_TA2_IO_012,
    output wire        mb1_FA1_TA1_IO_013_mb1_FB1_TA2_IO_013,
    output wire        mb1_FA1_TA1_IO_014_mb1_FB1_TA2_IO_016,
    output wire        mb1_FA1_TA1_IO_015_mb1_FB1_TA2_IO_017,
    output wire        mb1_FA1_TA1_IO_016_mb1_FB1_TA2_IO_014,
    output wire        mb1_FA1_TA1_IO_017_mb1_FB1_TA2_IO_015,
    output wire        mb1_FA1_TA1_IO_018_mb1_FB1_TA2_IO_032,
    output wire        mb1_FA1_TA1_IO_019_mb1_FB1_TA2_IO_033,
    output wire        mb1_FA1_TA1_IO_020_mb1_FB1_TA2_IO_030,
    output wire        mb1_FA1_TA1_IO_021_mb1_FB1_TA2_IO_031,
    output wire        mb1_FA1_TA1_IO_022_mb1_FB1_TA2_IO_008,
    output wire        mb1_FA1_TA1_IO_023_mb1_FB1_TA2_IO_009,
    output wire        mb1_FA1_TA1_IO_024_mb1_FB1_TA2_IO_026,
    output wire        mb1_FA1_TA1_IO_025_mb1_FB1_TA2_IO_027,
    output wire        mb1_FA1_TA1_IO_026_mb1_FB1_TA2_IO_024,
    output wire        mb1_FA1_TA1_IO_027_mb1_FB1_TA2_IO_025,
    output wire        mb1_FA1_TA1_IO_028_mb1_FB1_TA2_IO_042,
    output wire        mb1_FA1_TA1_IO_029_mb1_FB1_TA2_IO_043,
    output wire        mb1_FA1_TA1_IO_030_mb1_FB1_TA2_IO_020,
    output wire        mb1_FA1_TA1_IO_031_mb1_FB1_TA2_IO_021,
    output wire        mb1_FA1_TA1_IO_032_mb1_FB1_TA2_IO_018,
    output wire        mb1_FA1_TA1_IO_033_mb1_FB1_TA2_IO_019,
    output wire        mb1_FA1_TA1_IO_034_mb1_FB1_TA2_IO_036,
    output wire        mb1_FA1_TA1_IO_035_mb1_FB1_TA2_IO_037,
    output wire        mb1_FA1_TA1_IO_036_mb1_FB1_TA2_IO_034,
    output wire        mb1_FA1_TA1_IO_037_mb1_FB1_TA2_IO_035,
    output wire        mb1_FA1_TA1_IO_038_mb1_FB1_TA2_IO_052,
    output wire        mb1_FA1_TA1_IO_039_mb1_FB1_TA2_IO_053,
    output wire        mb1_FA1_TA1_IO_040_mb1_FB1_TA2_IO_050,
    output wire        mb1_FA1_TA1_IO_041_mb1_FB1_TA2_IO_051,
    output wire        mb1_FA1_TA1_IO_042_mb1_FB1_TA2_IO_028,
    output wire        mb1_FA1_TA1_IO_043_mb1_FB1_TA2_IO_029,
    output wire        mb1_FA1_TA1_IO_044_mb1_FB1_TA2_IO_046,
    output wire        mb1_FA1_TA1_IO_045_mb1_FB1_TA2_IO_047,
    output wire        mb1_FA1_TA1_IO_046_mb1_FB1_TA2_IO_044,
    output wire        mb1_FA1_TA1_IO_047_mb1_FB1_TA2_IO_045,
    output wire        mb1_FA1_TA1_IO_048_mb1_FB1_TA2_IO_062,
    output wire        mb1_FA1_TA1_IO_049_mb1_FB1_TA2_IO_063,
    output wire        mb1_FA1_TA1_IO_050_mb1_FB1_TA2_IO_040,
    output wire        mb1_FA1_TA1_IO_051_mb1_FB1_TA2_IO_041,
    output wire        mb1_FA1_TA1_IO_052_mb1_FB1_TA2_IO_038,
    output wire        mb1_FA1_TA1_IO_053_mb1_FB1_TA2_IO_039,
    output wire        mb1_FA1_TA1_IO_054_mb1_FB1_TA2_IO_056,
    output wire        mb1_FA1_TA1_IO_055_mb1_FB1_TA2_IO_057,
    output wire        mb1_FA1_TA1_IO_056_mb1_FB1_TA2_IO_054,
    output wire        mb1_FA1_TA1_IO_057_mb1_FB1_TA2_IO_055,
    output wire        mb1_FA1_TA1_IO_058_mb1_FB1_TA2_IO_072,
    output wire        mb1_FA1_TA1_IO_059_mb1_FB1_TA2_IO_073,
    output wire        mb1_FA1_TA1_IO_060_mb1_FB1_TA2_IO_070,
    output wire        mb1_FA1_TA1_IO_061_mb1_FB1_TA2_IO_071,
    output wire        mb1_FA1_TA1_IO_062_mb1_FB1_TA2_IO_048,
    output wire        mb1_FA1_TA1_IO_063_mb1_FB1_TA2_IO_049,
    output wire        mb1_FA1_TA1_IO_064_mb1_FB1_TA2_IO_066,
    output wire        mb1_FA1_TA1_IO_065_mb1_FB1_TA2_IO_067,
    output wire        mb1_FA1_TA1_IO_066_mb1_FB1_TA2_IO_064,
    output wire        mb1_FA1_TA1_IO_067_mb1_FB1_TA2_IO_065,
    output wire        mb1_FA1_TA1_IO_068_mb1_FB1_TA2_IO_082,
    output wire        mb1_FA1_TA1_IO_069_mb1_FB1_TA2_IO_083,
    output wire        mb1_FA1_TA1_IO_070_mb1_FB1_TA2_IO_060,
    output wire        mb1_FA1_TA1_IO_071_mb1_FB1_TA2_IO_061,
    output wire        mb1_FA1_TA1_IO_072_mb1_FB1_TA2_IO_058,
    output wire        mb1_FA1_TA1_IO_073_mb1_FB1_TA2_IO_059,
    output wire        mb1_FA1_TA1_IO_074_mb1_FB1_TA2_IO_076,
    output wire        mb1_FA1_TA1_IO_075_mb1_FB1_TA2_IO_077,
    output wire        mb1_FA1_TA1_IO_076_mb1_FB1_TA2_IO_074,
    output wire        mb1_FA1_TA1_IO_077_mb1_FB1_TA2_IO_075,
    output wire        mb1_FA1_TA1_IO_078_mb1_FB1_TA2_IO_092,
    output wire        mb1_FA1_TA1_IO_079_mb1_FB1_TA2_IO_093,
    output wire        mb1_FA1_TA1_IO_080_mb1_FB1_TA2_IO_090,
    output wire        mb1_FA1_TA1_IO_081_mb1_FB1_TA2_IO_091,
    output wire        mb1_FA1_TA1_IO_082_mb1_FB1_TA2_IO_068,
    output wire        mb1_FA1_TA1_IO_083_mb1_FB1_TA2_IO_069,
    output wire        mb1_FA1_TA1_IO_084_mb1_FB1_TA2_IO_086,
    output wire        mb1_FA1_TA1_IO_085_mb1_FB1_TA2_IO_087,
    output wire        mb1_FA1_TA1_IO_086_mb1_FB1_TA2_IO_084,
    output wire        mb1_FA1_TA1_IO_087_mb1_FB1_TA2_IO_085,
    output wire        mb1_FA1_TA1_IO_088_mb1_FB1_TA2_IO_102,
    output wire        mb1_FA1_TA1_IO_089_mb1_FB1_TA2_IO_103,
    output wire        mb1_FA1_TA1_IO_090_mb1_FB1_TA2_IO_080,
    output wire        mb1_FA1_TA1_IO_091_mb1_FB1_TA2_IO_081,
    output wire        mb1_FA1_TA1_IO_092_mb1_FB1_TA2_IO_078,
    output wire        mb1_FA1_TA1_IO_093_mb1_FB1_TA2_IO_079,
    output wire        mb1_FA1_TA1_IO_094_mb1_FB1_TA2_IO_096,
    output wire        mb1_FA1_TA1_IO_095_mb1_FB1_TA2_IO_097,
    output wire        mb1_FA1_TA1_IO_096_mb1_FB1_TA2_IO_094,
    output wire        mb1_FA1_TA1_IO_097_mb1_FB1_TA2_IO_095,
    output wire        mb1_FA1_TA1_IO_098_mb1_FB1_TA2_IO_112,
    output wire        mb1_FA1_TA1_IO_099_mb1_FB1_TA2_IO_113,
    output wire        mb1_FA1_TA1_IO_100_mb1_FB1_TA2_IO_110,
    output wire        mb1_FA1_TA1_IO_101_mb1_FB1_TA2_IO_111,
    output wire        mb1_FA1_TA1_IO_102_mb1_FB1_TA2_IO_088,
    output wire        mb1_FA1_TA1_IO_103_mb1_FB1_TA2_IO_089,
    output wire        mb1_FA1_TA1_IO_104_mb1_FB1_TA2_IO_106,
    output wire        mb1_FA1_TA1_IO_105_mb1_FB1_TA2_IO_107,
    output wire        mb1_FA1_TA1_IO_106_mb1_FB1_TA2_IO_104,
    output wire        mb1_FA1_TA1_IO_107_mb1_FB1_TA2_IO_105,
    output wire        mb1_FA1_TA1_IO_108_mb1_FB1_TA2_IO_122,
    output wire        mb1_FA1_TA1_IO_109_mb1_FB1_TA2_IO_123,
    output wire        mb1_FA1_TA1_IO_110_mb1_FB1_TA2_IO_100,
    output wire        mb1_FA1_TA1_IO_111_mb1_FB1_TA2_IO_101,
    output wire        mb1_FA1_TA1_IO_112_mb1_FB1_TA2_IO_098,
    output wire        mb1_FA1_TA1_IO_113_mb1_FB1_TA2_IO_099,
    output wire        mb1_FA1_TA1_IO_114_mb1_FB1_TA2_IO_116,
    output wire        mb1_FA1_TA1_IO_115_mb1_FB1_TA2_IO_117,
    output wire        mb1_FA1_TA1_IO_116_mb1_FB1_TA2_IO_114,
    output wire        mb1_FA1_TA1_IO_117_mb1_FB1_TA2_IO_115,
    output wire        mb1_FA1_TA1_IO_118_mb1_FB1_TA2_IO_132,
    output wire        mb1_FA1_TA1_IO_119_mb1_FB1_TA2_IO_133,
    output wire        mb1_FA1_TA1_IO_120_mb1_FB1_TA2_IO_130,
    output wire        mb1_FA1_TA1_IO_121_mb1_FB1_TA2_IO_131,
    output wire        mb1_FA1_TA1_IO_122_mb1_FB1_TA2_IO_108,
    output wire        mb1_FA1_TA1_IO_123_mb1_FB1_TA2_IO_109,
    output wire        mb1_FA1_TA1_IO_124_mb1_FB1_TA2_IO_126,
    output wire        mb1_FA1_TA1_IO_125_mb1_FB1_TA2_IO_127,
    output wire        mb1_FA1_TA1_IO_126_mb1_FB1_TA2_IO_124,
    output wire        mb1_FA1_TA1_IO_127_mb1_FB1_TA2_IO_125,
    output wire        mb1_FA1_TA1_IO_130_mb1_FB1_TA2_IO_120,
    output wire        mb1_FA1_TA1_IO_131_mb1_FB1_TA2_IO_121,
    output wire        mb1_FA1_TA1_IO_132_mb1_FB1_TA2_IO_118,
    output wire        mb1_FA1_TA1_IO_133_mb1_FB1_TA2_IO_119,
    output wire        mb1_FA1_TA1_IO_134_mb1_FB1_TA2_IO_136,
    output wire        mb1_FA1_TA1_IO_136_mb1_FB1_TA2_IO_134,
    output wire        mb1_FA1_TB0_CLKIO_N_0_mb1_FB1_TB2_CLKIO_N_7,
    output wire        mb1_FA1_TB0_CLKIO_N_1_mb1_FB1_TB2_CLKIO_N_6,
    output wire        mb1_FA1_TB0_CLKIO_N_2_mb1_FB1_TB2_CLKIO_N_4,
    output wire        mb1_FA1_TB0_CLKIO_N_3_mb1_FB1_TB2_CLKIO_N_3,
    output wire        mb1_FA1_TB0_CLKIO_N_4_mb1_FB1_TB2_CLKIO_N_2,
    output wire        mb1_FA1_TB0_CLKIO_N_5_mb1_FB1_TB2_IO_010,
    output wire        mb1_FA1_TB0_CLKIO_N_6_mb1_FB1_TB2_CLKIO_N_1,
    output wire        mb1_FA1_TB0_CLKIO_N_7_mb1_FB1_TB2_CLKIO_N_0,
    output wire        mb1_FA1_TB0_CLKIO_P_0_mb1_FB1_TB2_CLKIO_P_7,
    output wire        mb1_FA1_TB0_CLKIO_P_1_mb1_FB1_TB2_CLKIO_P_6,
    output wire        mb1_FA1_TB0_CLKIO_P_2_mb1_FB1_TB2_CLKIO_P_4,
    output wire        mb1_FA1_TB0_CLKIO_P_3_mb1_FB1_TB2_CLKIO_P_3,
    output wire        mb1_FA1_TB0_CLKIO_P_4_mb1_FB1_TB2_CLKIO_P_2,
    output wire        mb1_FA1_TB0_CLKIO_P_5_mb1_FB1_TB2_IO_011,
    output wire        mb1_FA1_TB0_CLKIO_P_6_mb1_FB1_TB2_CLKIO_P_1,
    output wire        mb1_FA1_TB0_CLKIO_P_7_mb1_FB1_TB2_CLKIO_P_0,
    output wire        mb1_FA1_TB0_IO_004_mb1_FB1_TB2_IO_006,
    output wire        mb1_FA1_TB0_IO_005_mb1_FB1_TB2_IO_007,
    output wire        mb1_FA1_TB0_IO_006_mb1_FB1_TB2_IO_004,
    output wire        mb1_FA1_TB0_IO_007_mb1_FB1_TB2_IO_005,
    output wire        mb1_FA1_TB0_IO_008_mb1_FB1_TB2_IO_022,
    output wire        mb1_FA1_TB0_IO_009_mb1_FB1_TB2_IO_023,
    output wire        mb1_FA1_TB0_IO_010_mb1_FB1_TB2_CLKIO_N_5,
    output wire        mb1_FA1_TB0_IO_011_mb1_FB1_TB2_CLKIO_P_5,
    output wire        mb1_FA1_TB0_IO_012_mb1_FB1_TB2_IO_012,
    output wire        mb1_FA1_TB0_IO_013_mb1_FB1_TB2_IO_013,
    output wire        mb1_FA1_TB0_IO_014_mb1_FB1_TB2_IO_016,
    output wire        mb1_FA1_TB0_IO_015_mb1_FB1_TB2_IO_017,
    output wire        mb1_FA1_TB0_IO_016_mb1_FB1_TB2_IO_014,
    output wire        mb1_FA1_TB0_IO_017_mb1_FB1_TB2_IO_015,
    output wire        mb1_FA1_TB0_IO_018_mb1_FB1_TB2_IO_032,
    output wire        mb1_FA1_TB0_IO_019_mb1_FB1_TB2_IO_033,
    output wire        mb1_FA1_TB0_IO_020_mb1_FB1_TB2_IO_030,
    output wire        mb1_FA1_TB0_IO_021_mb1_FB1_TB2_IO_031,
    output wire        mb1_FA1_TB0_IO_022_mb1_FB1_TB2_IO_008,
    output wire        mb1_FA1_TB0_IO_023_mb1_FB1_TB2_IO_009,
    output wire        mb1_FA1_TB0_IO_024_mb1_FB1_TB2_IO_026,
    output wire        mb1_FA1_TB0_IO_025_mb1_FB1_TB2_IO_027,
    output wire        mb1_FA1_TB0_IO_026_mb1_FB1_TB2_IO_024,
    output wire        mb1_FA1_TB0_IO_027_mb1_FB1_TB2_IO_025,
    output wire        mb1_FA1_TB0_IO_028_mb1_FB1_TB2_IO_042,
    output wire        mb1_FA1_TB0_IO_029_mb1_FB1_TB2_IO_043,
    output wire        mb1_FA1_TB0_IO_030_mb1_FB1_TB2_IO_020,
    output wire        mb1_FA1_TB0_IO_031_mb1_FB1_TB2_IO_021,
    output wire        mb1_FA1_TB0_IO_032_mb1_FB1_TB2_IO_018,
    output wire        mb1_FA1_TB0_IO_033_mb1_FB1_TB2_IO_019,
    output wire        mb1_FA1_TB0_IO_034_mb1_FB1_TB2_IO_036,
    output wire        mb1_FA1_TB0_IO_035_mb1_FB1_TB2_IO_037,
    output wire        mb1_FA1_TB0_IO_036_mb1_FB1_TB2_IO_034,
    output wire        mb1_FA1_TB0_IO_037_mb1_FB1_TB2_IO_035,
    output wire        mb1_FA1_TB0_IO_038_mb1_FB1_TB2_IO_052,
    output wire        mb1_FA1_TB0_IO_039_mb1_FB1_TB2_IO_053,
    output wire        mb1_FA1_TB0_IO_040_mb1_FB1_TB2_IO_050,
    output wire        mb1_FA1_TB0_IO_041_mb1_FB1_TB2_IO_051,
    output wire        mb1_FA1_TB0_IO_042_mb1_FB1_TB2_IO_028,
    output wire        mb1_FA1_TB0_IO_043_mb1_FB1_TB2_IO_029,
    output wire        mb1_FA1_TB0_IO_044_mb1_FB1_TB2_IO_046,
    output wire        mb1_FA1_TB0_IO_045_mb1_FB1_TB2_IO_047,
    output wire        mb1_FA1_TB0_IO_046_mb1_FB1_TB2_IO_044,
    output wire        mb1_FA1_TB0_IO_047_mb1_FB1_TB2_IO_045,
    output wire        mb1_FA1_TB0_IO_048_mb1_FB1_TB2_IO_062,
    output wire        mb1_FA1_TB0_IO_049_mb1_FB1_TB2_IO_063,
    output wire        mb1_FA1_TB0_IO_050_mb1_FB1_TB2_IO_040,
    output wire        mb1_FA1_TB0_IO_051_mb1_FB1_TB2_IO_041,
    output wire        mb1_FA1_TB0_IO_052_mb1_FB1_TB2_IO_038,
    output wire        mb1_FA1_TB0_IO_053_mb1_FB1_TB2_IO_039,
    output wire        mb1_FA1_TB0_IO_054_mb1_FB1_TB2_IO_056,
    output wire        mb1_FA1_TB0_IO_055_mb1_FB1_TB2_IO_057,
    output wire        mb1_FA1_TB0_IO_056_mb1_FB1_TB2_IO_054,
    output wire        mb1_FA1_TB0_IO_057_mb1_FB1_TB2_IO_055,
    output wire        mb1_FA1_TB0_IO_058_mb1_FB1_TB2_IO_072,
    output wire        mb1_FA1_TB0_IO_059_mb1_FB1_TB2_IO_073,
    output wire        mb1_FA1_TB0_IO_060_mb1_FB1_TB2_IO_070,
    output wire        mb1_FA1_TB0_IO_061_mb1_FB1_TB2_IO_071,
    output wire        mb1_FA1_TB0_IO_062_mb1_FB1_TB2_IO_048,
    output wire        mb1_FA1_TB0_IO_063_mb1_FB1_TB2_IO_049,
    output wire        mb1_FA1_TB0_IO_064_mb1_FB1_TB2_IO_066,
    output wire        mb1_FA1_TB0_IO_065_mb1_FB1_TB2_IO_067,
    output wire        mb1_FA1_TB0_IO_066_mb1_FB1_TB2_IO_064,
    output wire        mb1_FA1_TB0_IO_067_mb1_FB1_TB2_IO_065,
    output wire        mb1_FA1_TB0_IO_068_mb1_FB1_TB2_IO_082,
    output wire        mb1_FA1_TB0_IO_069_mb1_FB1_TB2_IO_083,
    output wire        mb1_FA1_TB0_IO_070_mb1_FB1_TB2_IO_060,
    output wire        mb1_FA1_TB0_IO_071_mb1_FB1_TB2_IO_061,
    output wire        mb1_FA1_TB0_IO_072_mb1_FB1_TB2_IO_058,
    output wire        mb1_FA1_TB0_IO_073_mb1_FB1_TB2_IO_059,
    output wire        mb1_FA1_TB0_IO_074_mb1_FB1_TB2_IO_076,
    output wire        mb1_FA1_TB0_IO_075_mb1_FB1_TB2_IO_077,
    output wire        mb1_FA1_TB0_IO_076_mb1_FB1_TB2_IO_074,
    output wire        mb1_FA1_TB0_IO_077_mb1_FB1_TB2_IO_075,
    output wire        mb1_FA1_TB0_IO_078_mb1_FB1_TB2_IO_092,
    output wire        mb1_FA1_TB0_IO_079_mb1_FB1_TB2_IO_093,
    output wire        mb1_FA1_TB0_IO_080_mb1_FB1_TB2_IO_090,
    output wire        mb1_FA1_TB0_IO_081_mb1_FB1_TB2_IO_091,
    output wire        mb1_FA1_TB0_IO_082_mb1_FB1_TB2_IO_068,
    output wire        mb1_FA1_TB0_IO_083_mb1_FB1_TB2_IO_069,
    output wire        mb1_FA1_TB0_IO_084_mb1_FB1_TB2_IO_086,
    output wire        mb1_FA1_TB0_IO_085_mb1_FB1_TB2_IO_087,
    output wire        mb1_FA1_TB0_IO_086_mb1_FB1_TB2_IO_084,
    output wire        mb1_FA1_TB0_IO_087_mb1_FB1_TB2_IO_085,
    output wire        mb1_FA1_TB0_IO_088_mb1_FB1_TB2_IO_102,
    output wire        mb1_FA1_TB0_IO_089_mb1_FB1_TB2_IO_103,
    output wire        mb1_FA1_TB0_IO_090_mb1_FB1_TB2_IO_080,
    output wire        mb1_FA1_TB0_IO_091_mb1_FB1_TB2_IO_081,
    output wire        mb1_FA1_TB0_IO_092_mb1_FB1_TB2_IO_078,
    output wire        mb1_FA1_TB0_IO_093_mb1_FB1_TB2_IO_079,
    output wire        mb1_FA1_TB0_IO_094_mb1_FB1_TB2_IO_096,
    output wire        mb1_FA1_TB0_IO_095_mb1_FB1_TB2_IO_097,
    output wire        mb1_FA1_TB0_IO_096_mb1_FB1_TB2_IO_094,
    output wire        mb1_FA1_TB0_IO_097_mb1_FB1_TB2_IO_095,
    output wire        mb1_FA1_TB0_IO_098_mb1_FB1_TB2_IO_112,
    output wire        mb1_FA1_TB0_IO_099_mb1_FB1_TB2_IO_113,
    output wire        mb1_FA1_TB0_IO_100_mb1_FB1_TB2_IO_110,
    output wire        mb1_FA1_TB0_IO_101_mb1_FB1_TB2_IO_111,
    output wire        mb1_FA1_TB0_IO_102_mb1_FB1_TB2_IO_088,
    output wire        mb1_FA1_TB0_IO_103_mb1_FB1_TB2_IO_089,
    output wire        mb1_FA1_TB0_IO_104_mb1_FB1_TB2_IO_106,
    output wire        mb1_FA1_TB0_IO_105_mb1_FB1_TB2_IO_107,
    output wire        mb1_FA1_TB0_IO_106_mb1_FB1_TB2_IO_104,
    output wire        mb1_FA1_TB0_IO_107_mb1_FB1_TB2_IO_105,
    output wire        mb1_FA1_TB0_IO_108_mb1_FB1_TB2_IO_122,
    output wire        mb1_FA1_TB0_IO_109_mb1_FB1_TB2_IO_123,
    output wire        mb1_FA1_TB0_IO_110_mb1_FB1_TB2_IO_100,
    output wire        mb1_FA1_TB0_IO_111_mb1_FB1_TB2_IO_101,
    output wire        mb1_FA1_TB0_IO_112_mb1_FB1_TB2_IO_098,
    output wire        mb1_FA1_TB0_IO_113_mb1_FB1_TB2_IO_099,
    output wire        mb1_FA1_TB0_IO_114_mb1_FB1_TB2_IO_116,
    output wire        mb1_FA1_TB0_IO_115_mb1_FB1_TB2_IO_117,
    output wire        mb1_FA1_TB0_IO_116_mb1_FB1_TB2_IO_114,
    output wire        mb1_FA1_TB0_IO_117_mb1_FB1_TB2_IO_115,
    output wire        mb1_FA1_TB0_IO_118_mb1_FB1_TB2_IO_132,
    output wire        mb1_FA1_TB0_IO_119_mb1_FB1_TB2_IO_133,
    output wire        mb1_FA1_TB0_IO_120_mb1_FB1_TB2_IO_130,
    output wire        mb1_FA1_TB0_IO_121_mb1_FB1_TB2_IO_131,
    output wire        mb1_FA1_TB0_IO_122_mb1_FB1_TB2_IO_108,
    output wire        mb1_FA1_TB0_IO_123_mb1_FB1_TB2_IO_109,
    output wire        mb1_FA1_TB0_IO_124_mb1_FB1_TB2_IO_126,
    output wire        mb1_FA1_TB0_IO_125_mb1_FB1_TB2_IO_127,
    output wire        mb1_FA1_TB0_IO_126_mb1_FB1_TB2_IO_124,
    output wire        mb1_FA1_TB0_IO_127_mb1_FB1_TB2_IO_125,
    output wire        mb1_FA1_TB0_IO_130_mb1_FB1_TB2_IO_120,
    output wire        mb1_FA1_TB0_IO_131_mb1_FB1_TB2_IO_121,
    output wire        mb1_FA1_TB0_IO_132_mb1_FB1_TB2_IO_118,
    output wire        mb1_FA1_TB0_IO_133_mb1_FB1_TB2_IO_119,
    output wire        mb1_FA1_TB0_IO_134_mb1_FB1_TB2_IO_136,
    output wire        mb1_FA1_TB0_IO_136_mb1_FB1_TB2_IO_134,
    output wire        mb1_FA1_TB1_CLKIO_N_0_mb1_FB1_BB1_CLKIO_N_7,
    output wire        mb1_FA1_TB1_CLKIO_N_1_mb1_FB1_BB1_CLKIO_N_6,
    output wire        mb1_FA1_TB1_CLKIO_N_2_mb1_FB1_BB1_CLKIO_N_4,
    output wire        mb1_FA1_TB1_CLKIO_N_3_mb1_FB1_BB1_CLKIO_N_3,
    output wire        mb1_FA1_TB1_CLKIO_N_4_mb1_FB1_BB1_CLKIO_N_2,
    output wire        mb1_FA1_TB1_CLKIO_N_5_mb1_FB1_BB1_IO_010,
    output wire        mb1_FA1_TB1_CLKIO_N_6_mb1_FB1_BB1_CLKIO_N_1,
    output wire        mb1_FA1_TB1_CLKIO_N_7_mb1_FB1_BB1_CLKIO_N_0,
    output wire        mb1_FA1_TB1_CLKIO_P_0_mb1_FB1_BB1_CLKIO_P_7,
    output wire        mb1_FA1_TB1_CLKIO_P_1_mb1_FB1_BB1_CLKIO_P_6,
    output wire        mb1_FA1_TB1_CLKIO_P_2_mb1_FB1_BB1_CLKIO_P_4,
    output wire        mb1_FA1_TB1_CLKIO_P_3_mb1_FB1_BB1_CLKIO_P_3,
    output wire        mb1_FA1_TB1_CLKIO_P_4_mb1_FB1_BB1_CLKIO_P_2,
    output wire        mb1_FA1_TB1_CLKIO_P_5_mb1_FB1_BB1_IO_011,
    output wire        mb1_FA1_TB1_CLKIO_P_6_mb1_FB1_BB1_CLKIO_P_1,
    output wire        mb1_FA1_TB1_CLKIO_P_7_mb1_FB1_BB1_CLKIO_P_0,
    output wire        mb1_FA1_TB1_IO_004_mb1_FB1_BB1_IO_006,
    output wire        mb1_FA1_TB1_IO_005_mb1_FB1_BB1_IO_007,
    output wire        mb1_FA1_TB1_IO_006_mb1_FB1_BB1_IO_004,
    output wire        mb1_FA1_TB1_IO_007_mb1_FB1_BB1_IO_005,
    output wire        mb1_FA1_TB1_IO_008_mb1_FB1_BB1_IO_022,
    output wire        mb1_FA1_TB1_IO_009_mb1_FB1_BB1_IO_023,
    output wire        mb1_FA1_TB1_IO_010_mb1_FB1_BB1_CLKIO_N_5,
    output wire        mb1_FA1_TB1_IO_011_mb1_FB1_BB1_CLKIO_P_5,
    output wire        mb1_FA1_TB1_IO_012_mb1_FB1_BB1_IO_012,
    output wire        mb1_FA1_TB1_IO_013_mb1_FB1_BB1_IO_013,
    output wire        mb1_FA1_TB1_IO_014_mb1_FB1_BB1_IO_016,
    output wire        mb1_FA1_TB1_IO_015_mb1_FB1_BB1_IO_017,
    output wire        mb1_FA1_TB1_IO_016_mb1_FB1_BB1_IO_014,
    output wire        mb1_FA1_TB1_IO_017_mb1_FB1_BB1_IO_015,
    output wire        mb1_FA1_TB1_IO_018_mb1_FB1_BB1_IO_032,
    output wire        mb1_FA1_TB1_IO_019_mb1_FB1_BB1_IO_033,
    output wire        mb1_FA1_TB1_IO_020_mb1_FB1_BB1_IO_030,
    output wire        mb1_FA1_TB1_IO_021_mb1_FB1_BB1_IO_031,
    output wire        mb1_FA1_TB1_IO_022_mb1_FB1_BB1_IO_008,
    output wire        mb1_FA1_TB1_IO_023_mb1_FB1_BB1_IO_009,
    output wire        mb1_FA1_TB1_IO_024_mb1_FB1_BB1_IO_026,
    output wire        mb1_FA1_TB1_IO_025_mb1_FB1_BB1_IO_027,
    output wire        mb1_FA1_TB1_IO_026_mb1_FB1_BB1_IO_024,
    output wire        mb1_FA1_TB1_IO_027_mb1_FB1_BB1_IO_025,
    output wire        mb1_FA1_TB1_IO_028_mb1_FB1_BB1_IO_042,
    output wire        mb1_FA1_TB1_IO_029_mb1_FB1_BB1_IO_043,
    output wire        mb1_FA1_TB1_IO_030_mb1_FB1_BB1_IO_020,
    output wire        mb1_FA1_TB1_IO_031_mb1_FB1_BB1_IO_021,
    output wire        mb1_FA1_TB1_IO_032_mb1_FB1_BB1_IO_018,
    output wire        mb1_FA1_TB1_IO_033_mb1_FB1_BB1_IO_019,
    output wire        mb1_FA1_TB1_IO_034_mb1_FB1_BB1_IO_036,
    output wire        mb1_FA1_TB1_IO_035_mb1_FB1_BB1_IO_037,
    output wire        mb1_FA1_TB1_IO_036_mb1_FB1_BB1_IO_034,
    output wire        mb1_FA1_TB1_IO_037_mb1_FB1_BB1_IO_035,
    output wire        mb1_FA1_TB1_IO_038_mb1_FB1_BB1_IO_052,
    output wire        mb1_FA1_TB1_IO_039_mb1_FB1_BB1_IO_053,
    output wire        mb1_FA1_TB1_IO_040_mb1_FB1_BB1_IO_050,
    output wire        mb1_FA1_TB1_IO_041_mb1_FB1_BB1_IO_051,
    output wire        mb1_FA1_TB1_IO_042_mb1_FB1_BB1_IO_028,
    output wire        mb1_FA1_TB1_IO_043_mb1_FB1_BB1_IO_029,
    output wire        mb1_FA1_TB1_IO_044_mb1_FB1_BB1_IO_046,
    output wire        mb1_FA1_TB1_IO_045_mb1_FB1_BB1_IO_047,
    output wire        mb1_FA1_TB1_IO_046_mb1_FB1_BB1_IO_044,
    output wire        mb1_FA1_TB1_IO_047_mb1_FB1_BB1_IO_045,
    output wire        mb1_FA1_TB1_IO_048_mb1_FB1_BB1_IO_062,
    output wire        mb1_FA1_TB1_IO_049_mb1_FB1_BB1_IO_063,
    output wire        mb1_FA1_TB1_IO_050_mb1_FB1_BB1_IO_040,
    output wire        mb1_FA1_TB1_IO_051_mb1_FB1_BB1_IO_041,
    output wire        mb1_FA1_TB1_IO_052_mb1_FB1_BB1_IO_038,
    output wire        mb1_FA1_TB1_IO_053_mb1_FB1_BB1_IO_039,
    output wire        mb1_FA1_TB1_IO_054_mb1_FB1_BB1_IO_056,
    output wire        mb1_FA1_TB1_IO_055_mb1_FB1_BB1_IO_057,
    output wire        mb1_FA1_TB1_IO_056_mb1_FB1_BB1_IO_054,
    output wire        mb1_FA1_TB1_IO_057_mb1_FB1_BB1_IO_055,
    output wire        mb1_FA1_TB1_IO_058_mb1_FB1_BB1_IO_072,
    output wire        mb1_FA1_TB1_IO_059_mb1_FB1_BB1_IO_073,
    output wire        mb1_FA1_TB1_IO_060_mb1_FB1_BB1_IO_070,
    output wire        mb1_FA1_TB1_IO_061_mb1_FB1_BB1_IO_071,
    output wire        mb1_FA1_TB1_IO_062_mb1_FB1_BB1_IO_048,
    output wire        mb1_FA1_TB1_IO_063_mb1_FB1_BB1_IO_049,
    output wire        mb1_FA1_TB1_IO_064_mb1_FB1_BB1_IO_066,
    output wire        mb1_FA1_TB1_IO_065_mb1_FB1_BB1_IO_067,
    output wire        mb1_FA1_TB1_IO_066_mb1_FB1_BB1_IO_064,
    output wire        mb1_FA1_TB1_IO_067_mb1_FB1_BB1_IO_065,
    output wire        mb1_FA1_TB1_IO_068_mb1_FB1_BB1_IO_082,
    output wire        mb1_FA1_TB1_IO_069_mb1_FB1_BB1_IO_083,
    output wire        mb1_FA1_TB1_IO_070_mb1_FB1_BB1_IO_060,
    output wire        mb1_FA1_TB1_IO_071_mb1_FB1_BB1_IO_061,
    output wire        mb1_FA1_TB1_IO_072_mb1_FB1_BB1_IO_058,
    output wire        mb1_FA1_TB1_IO_073_mb1_FB1_BB1_IO_059,
    output wire        mb1_FA1_TB1_IO_074_mb1_FB1_BB1_IO_076,
    output wire        mb1_FA1_TB1_IO_075_mb1_FB1_BB1_IO_077,
    output wire        mb1_FA1_TB1_IO_076_mb1_FB1_BB1_IO_074,
    output wire        mb1_FA1_TB1_IO_077_mb1_FB1_BB1_IO_075,
    output wire        mb1_FA1_TB1_IO_078_mb1_FB1_BB1_IO_092,
    output wire        mb1_FA1_TB1_IO_079_mb1_FB1_BB1_IO_093,
    output wire        mb1_FA1_TB1_IO_080_mb1_FB1_BB1_IO_090,
    output wire        mb1_FA1_TB1_IO_081_mb1_FB1_BB1_IO_091,
    output wire        mb1_FA1_TB1_IO_082_mb1_FB1_BB1_IO_068,
    output wire        mb1_FA1_TB1_IO_083_mb1_FB1_BB1_IO_069,
    output wire        mb1_FA1_TB1_IO_084_mb1_FB1_BB1_IO_086,
    output wire        mb1_FA1_TB1_IO_085_mb1_FB1_BB1_IO_087,
    output wire        mb1_FA1_TB1_IO_086_mb1_FB1_BB1_IO_084,
    output wire        mb1_FA1_TB1_IO_087_mb1_FB1_BB1_IO_085,
    output wire        mb1_FA1_TB1_IO_088_mb1_FB1_BB1_IO_102,
    output wire        mb1_FA1_TB1_IO_089_mb1_FB1_BB1_IO_103,
    output wire        mb1_FA1_TB1_IO_090_mb1_FB1_BB1_IO_080,
    output wire        mb1_FA1_TB1_IO_091_mb1_FB1_BB1_IO_081,
    output wire        mb1_FA1_TB1_IO_092_mb1_FB1_BB1_IO_078,
    output wire        mb1_FA1_TB1_IO_093_mb1_FB1_BB1_IO_079,
    output wire        mb1_FA1_TB1_IO_094_mb1_FB1_BB1_IO_096,
    output wire        mb1_FA1_TB1_IO_095_mb1_FB1_BB1_IO_097,
    output wire        mb1_FA1_TB1_IO_096_mb1_FB1_BB1_IO_094,
    output wire        mb1_FA1_TB1_IO_097_mb1_FB1_BB1_IO_095,
    output wire        mb1_FA1_TB1_IO_098_mb1_FB1_BB1_IO_112,
    output wire        mb1_FA1_TB1_IO_099_mb1_FB1_BB1_IO_113,
    output wire        mb1_FA1_TB1_IO_100_mb1_FB1_BB1_IO_110,
    output wire        mb1_FA1_TB1_IO_101_mb1_FB1_BB1_IO_111,
    output wire        mb1_FA1_TB1_IO_102_mb1_FB1_BB1_IO_088,
    output wire        mb1_FA1_TB1_IO_103_mb1_FB1_BB1_IO_089,
    output wire        mb1_FA1_TB1_IO_104_mb1_FB1_BB1_IO_106,
    output wire        mb1_FA1_TB1_IO_105_mb1_FB1_BB1_IO_107,
    output wire        mb1_FA1_TB1_IO_106_mb1_FB1_BB1_IO_104,
    output wire        mb1_FA1_TB1_IO_107_mb1_FB1_BB1_IO_105,
    output wire        mb1_FA1_TB1_IO_108_mb1_FB1_BB1_IO_122,
    output wire        mb1_FA1_TB1_IO_109_mb1_FB1_BB1_IO_123,
    output wire        mb1_FA1_TB1_IO_110_mb1_FB1_BB1_IO_100,
    output wire        mb1_FA1_TB1_IO_111_mb1_FB1_BB1_IO_101,
    output wire        mb1_FA1_TB1_IO_112_mb1_FB1_BB1_IO_098,
    output wire        mb1_FA1_TB1_IO_113_mb1_FB1_BB1_IO_099,
    output wire        mb1_FA1_TB1_IO_114_mb1_FB1_BB1_IO_116,
    output wire        mb1_FA1_TB1_IO_115_mb1_FB1_BB1_IO_117,
    output wire        mb1_FA1_TB1_IO_116_mb1_FB1_BB1_IO_114,
    output wire        mb1_FA1_TB1_IO_117_mb1_FB1_BB1_IO_115,
    output wire        mb1_FA1_TB1_IO_118_mb1_FB1_BB1_IO_132,
    output wire        mb1_FA1_TB1_IO_119_mb1_FB1_BB1_IO_133,
    output wire        mb1_FA1_TB1_IO_120_mb1_FB1_BB1_IO_130,
    output wire        mb1_FA1_TB1_IO_121_mb1_FB1_BB1_IO_131,
    output wire        mb1_FA1_TB1_IO_122_mb1_FB1_BB1_IO_108,
    output wire        mb1_FA1_TB1_IO_123_mb1_FB1_BB1_IO_109,
    output wire        mb1_FA1_TB1_IO_124_mb1_FB1_BB1_IO_126,
    output wire        mb1_FA1_TB1_IO_125_mb1_FB1_BB1_IO_127,
    output wire        mb1_FA1_TB1_IO_126_mb1_FB1_BB1_IO_124,
    output wire        mb1_FA1_TB1_IO_127_mb1_FB1_BB1_IO_125,
    output wire        mb1_FA1_TB1_IO_130_mb1_FB1_BB1_IO_120,
    output wire        mb1_FA1_TB1_IO_131_mb1_FB1_BB1_IO_121,
    output wire        mb1_FA1_TB1_IO_132_mb1_FB1_BB1_IO_118,
    output wire        mb1_FA1_TB1_IO_133_mb1_FB1_BB1_IO_119,
    output wire        mb1_FA1_TB1_IO_134_mb1_FB1_BB1_IO_136,
    output wire        mb1_FA1_TB1_IO_136_mb1_FB1_BB1_IO_134,
    output wire        mb1_FA1_TB2_CLKIO_N_0_mb1_FB2_BB1_CLKIO_N_7,
    output wire        mb1_FA1_TB2_CLKIO_N_1_mb1_FB2_BB1_CLKIO_N_6,
    output wire        mb1_FA1_TB2_CLKIO_N_2_mb1_FB2_BB1_CLKIO_N_4,
    output wire        mb1_FA1_TB2_CLKIO_N_3_mb1_FB2_BB1_CLKIO_N_3,
    output wire        mb1_FA1_TB2_CLKIO_N_4_mb1_FB2_BB1_CLKIO_N_2,
    output wire        mb1_FA1_TB2_CLKIO_N_5_mb1_FB2_BB1_IO_010,
    output wire        mb1_FA1_TB2_CLKIO_N_6_mb1_FB2_BB1_CLKIO_N_1,
    output wire        mb1_FA1_TB2_CLKIO_N_7_mb1_FB2_BB1_CLKIO_N_0,
    output wire        mb1_FA1_TB2_CLKIO_P_0_mb1_FB2_BB1_CLKIO_P_7,
    output wire        mb1_FA1_TB2_CLKIO_P_1_mb1_FB2_BB1_CLKIO_P_6,
    output wire        mb1_FA1_TB2_CLKIO_P_2_mb1_FB2_BB1_CLKIO_P_4,
    output wire        mb1_FA1_TB2_CLKIO_P_3_mb1_FB2_BB1_CLKIO_P_3,
    output wire        mb1_FA1_TB2_CLKIO_P_4_mb1_FB2_BB1_CLKIO_P_2,
    output wire        mb1_FA1_TB2_CLKIO_P_5_mb1_FB2_BB1_IO_011,
    output wire        mb1_FA1_TB2_CLKIO_P_6_mb1_FB2_BB1_CLKIO_P_1,
    output wire        mb1_FA1_TB2_CLKIO_P_7_mb1_FB2_BB1_CLKIO_P_0,
    output wire        mb1_FA1_TB2_IO_004_mb1_FB2_BB1_IO_006,
    output wire        mb1_FA1_TB2_IO_005_mb1_FB2_BB1_IO_007,
    output wire        mb1_FA1_TB2_IO_006_mb1_FB2_BB1_IO_004,
    output wire        mb1_FA1_TB2_IO_007_mb1_FB2_BB1_IO_005,
    output wire        mb1_FA1_TB2_IO_008_mb1_FB2_BB1_IO_022,
    output wire        mb1_FA1_TB2_IO_009_mb1_FB2_BB1_IO_023,
    output wire        mb1_FA1_TB2_IO_010_mb1_FB2_BB1_CLKIO_N_5,
    output wire        mb1_FA1_TB2_IO_011_mb1_FB2_BB1_CLKIO_P_5,
    output wire        mb1_FA1_TB2_IO_012_mb1_FB2_BB1_IO_012,
    output wire        mb1_FA1_TB2_IO_013_mb1_FB2_BB1_IO_013,
    output wire        mb1_FA1_TB2_IO_014_mb1_FB2_BB1_IO_016,
    output wire        mb1_FA1_TB2_IO_015_mb1_FB2_BB1_IO_017,
    output wire        mb1_FA1_TB2_IO_016_mb1_FB2_BB1_IO_014,
    output wire        mb1_FA1_TB2_IO_017_mb1_FB2_BB1_IO_015,
    output wire        mb1_FA1_TB2_IO_018_mb1_FB2_BB1_IO_032,
    output wire        mb1_FA1_TB2_IO_019_mb1_FB2_BB1_IO_033,
    output wire        mb1_FA1_TB2_IO_020_mb1_FB2_BB1_IO_030,
    output wire        mb1_FA1_TB2_IO_021_mb1_FB2_BB1_IO_031,
    output wire        mb1_FA1_TB2_IO_022_mb1_FB2_BB1_IO_008,
    output wire        mb1_FA1_TB2_IO_023_mb1_FB2_BB1_IO_009,
    output wire        mb1_FA1_TB2_IO_024_mb1_FB2_BB1_IO_026,
    output wire        mb1_FA1_TB2_IO_025_mb1_FB2_BB1_IO_027,
    output wire        mb1_FA1_TB2_IO_026_mb1_FB2_BB1_IO_024,
    output wire        mb1_FA1_TB2_IO_027_mb1_FB2_BB1_IO_025,
    output wire        mb1_FA1_TB2_IO_028_mb1_FB2_BB1_IO_042,
    output wire        mb1_FA1_TB2_IO_029_mb1_FB2_BB1_IO_043,
    output wire        mb1_FA1_TB2_IO_030_mb1_FB2_BB1_IO_020,
    output wire        mb1_FA1_TB2_IO_031_mb1_FB2_BB1_IO_021,
    output wire        mb1_FA1_TB2_IO_032_mb1_FB2_BB1_IO_018,
    output wire        mb1_FA1_TB2_IO_033_mb1_FB2_BB1_IO_019,
    output wire        mb1_FA1_TB2_IO_034_mb1_FB2_BB1_IO_036,
    output wire        mb1_FA1_TB2_IO_035_mb1_FB2_BB1_IO_037,
    output wire        mb1_FA1_TB2_IO_036_mb1_FB2_BB1_IO_034,
    output wire        mb1_FA1_TB2_IO_037_mb1_FB2_BB1_IO_035,
    output wire        mb1_FA1_TB2_IO_038_mb1_FB2_BB1_IO_052,
    output wire        mb1_FA1_TB2_IO_039_mb1_FB2_BB1_IO_053,
    output wire        mb1_FA1_TB2_IO_040_mb1_FB2_BB1_IO_050,
    output wire        mb1_FA1_TB2_IO_041_mb1_FB2_BB1_IO_051,
    output wire        mb1_FA1_TB2_IO_042_mb1_FB2_BB1_IO_028,
    output wire        mb1_FA1_TB2_IO_043_mb1_FB2_BB1_IO_029,
    output wire        mb1_FA1_TB2_IO_044_mb1_FB2_BB1_IO_046,
    output wire        mb1_FA1_TB2_IO_045_mb1_FB2_BB1_IO_047,
    output wire        mb1_FA1_TB2_IO_046_mb1_FB2_BB1_IO_044,
    output wire        mb1_FA1_TB2_IO_047_mb1_FB2_BB1_IO_045,
    output wire        mb1_FA1_TB2_IO_048_mb1_FB2_BB1_IO_062,
    output wire        mb1_FA1_TB2_IO_049_mb1_FB2_BB1_IO_063,
    output wire        mb1_FA1_TB2_IO_050_mb1_FB2_BB1_IO_040,
    output wire        mb1_FA1_TB2_IO_051_mb1_FB2_BB1_IO_041,
    output wire        mb1_FA1_TB2_IO_052_mb1_FB2_BB1_IO_038,
    output wire        mb1_FA1_TB2_IO_053_mb1_FB2_BB1_IO_039,
    output wire        mb1_FA1_TB2_IO_054_mb1_FB2_BB1_IO_056,
    output wire        mb1_FA1_TB2_IO_055_mb1_FB2_BB1_IO_057,
    output wire        mb1_FA1_TB2_IO_056_mb1_FB2_BB1_IO_054,
    output wire        mb1_FA1_TB2_IO_057_mb1_FB2_BB1_IO_055,
    output wire        mb1_FA1_TB2_IO_058_mb1_FB2_BB1_IO_072,
    output wire        mb1_FA1_TB2_IO_059_mb1_FB2_BB1_IO_073,
    output wire        mb1_FA1_TB2_IO_060_mb1_FB2_BB1_IO_070,
    output wire        mb1_FA1_TB2_IO_061_mb1_FB2_BB1_IO_071,
    output wire        mb1_FA1_TB2_IO_062_mb1_FB2_BB1_IO_048,
    output wire        mb1_FA1_TB2_IO_063_mb1_FB2_BB1_IO_049,
    output wire        mb1_FA1_TB2_IO_064_mb1_FB2_BB1_IO_066,
    output wire        mb1_FA1_TB2_IO_065_mb1_FB2_BB1_IO_067,
    output wire        mb1_FA1_TB2_IO_066_mb1_FB2_BB1_IO_064,
    output wire        mb1_FA1_TB2_IO_067_mb1_FB2_BB1_IO_065,
    output wire        mb1_FA1_TB2_IO_068_mb1_FB2_BB1_IO_082,
    output wire        mb1_FA1_TB2_IO_069_mb1_FB2_BB1_IO_083,
    output wire        mb1_FA1_TB2_IO_070_mb1_FB2_BB1_IO_060,
    output wire        mb1_FA1_TB2_IO_071_mb1_FB2_BB1_IO_061,
    output wire        mb1_FA1_TB2_IO_072_mb1_FB2_BB1_IO_058,
    output wire        mb1_FA1_TB2_IO_073_mb1_FB2_BB1_IO_059,
    output wire        mb1_FA1_TB2_IO_074_mb1_FB2_BB1_IO_076,
    output wire        mb1_FA1_TB2_IO_075_mb1_FB2_BB1_IO_077,
    output wire        mb1_FA1_TB2_IO_076_mb1_FB2_BB1_IO_074,
    output wire        mb1_FA1_TB2_IO_077_mb1_FB2_BB1_IO_075,
    output wire        mb1_FA1_TB2_IO_078_mb1_FB2_BB1_IO_092,
    output wire        mb1_FA1_TB2_IO_079_mb1_FB2_BB1_IO_093,
    output wire        mb1_FA1_TB2_IO_080_mb1_FB2_BB1_IO_090,
    output wire        mb1_FA1_TB2_IO_081_mb1_FB2_BB1_IO_091,
    output wire        mb1_FA1_TB2_IO_082_mb1_FB2_BB1_IO_068,
    output wire        mb1_FA1_TB2_IO_083_mb1_FB2_BB1_IO_069,
    output wire        mb1_FA1_TB2_IO_084_mb1_FB2_BB1_IO_086,
    output wire        mb1_FA1_TB2_IO_085_mb1_FB2_BB1_IO_087,
    output wire        mb1_FA1_TB2_IO_086_mb1_FB2_BB1_IO_084,
    output wire        mb1_FA1_TB2_IO_087_mb1_FB2_BB1_IO_085,
    output wire        mb1_FA1_TB2_IO_088_mb1_FB2_BB1_IO_102,
    output wire        mb1_FA1_TB2_IO_089_mb1_FB2_BB1_IO_103,
    output wire        mb1_FA1_TB2_IO_090_mb1_FB2_BB1_IO_080,
    output wire        mb1_FA1_TB2_IO_091_mb1_FB2_BB1_IO_081,
    output wire        mb1_FA1_TB2_IO_092_mb1_FB2_BB1_IO_078,
    output wire        mb1_FA1_TB2_IO_093_mb1_FB2_BB1_IO_079,
    output wire        mb1_FA1_TB2_IO_094_mb1_FB2_BB1_IO_096,
    output wire        mb1_FA1_TB2_IO_095_mb1_FB2_BB1_IO_097,
    output wire        mb1_FA1_TB2_IO_096_mb1_FB2_BB1_IO_094,
    output wire        mb1_FA1_TB2_IO_097_mb1_FB2_BB1_IO_095,
    output wire        mb1_FA1_TB2_IO_098_mb1_FB2_BB1_IO_112,
    output wire        mb1_FA1_TB2_IO_099_mb1_FB2_BB1_IO_113,
    output wire        mb1_FA1_TB2_IO_100_mb1_FB2_BB1_IO_110,
    output wire        mb1_FA1_TB2_IO_101_mb1_FB2_BB1_IO_111,
    output wire        mb1_FA1_TB2_IO_102_mb1_FB2_BB1_IO_088,
    output wire        mb1_FA1_TB2_IO_103_mb1_FB2_BB1_IO_089,
    output wire        mb1_FA1_TB2_IO_104_mb1_FB2_BB1_IO_106,
    output wire        mb1_FA1_TB2_IO_105_mb1_FB2_BB1_IO_107,
    output wire        mb1_FA1_TB2_IO_106_mb1_FB2_BB1_IO_104,
    output wire        mb1_FA1_TB2_IO_107_mb1_FB2_BB1_IO_105,
    output wire        mb1_FA1_TB2_IO_108_mb1_FB2_BB1_IO_122,
    output wire        mb1_FA1_TB2_IO_109_mb1_FB2_BB1_IO_123,
    output wire        mb1_FA1_TB2_IO_110_mb1_FB2_BB1_IO_100,
    output wire        mb1_FA1_TB2_IO_111_mb1_FB2_BB1_IO_101,
    output wire        mb1_FA1_TB2_IO_112_mb1_FB2_BB1_IO_098,
    output wire        mb1_FA1_TB2_IO_113_mb1_FB2_BB1_IO_099,
    output wire        mb1_FA1_TB2_IO_114_mb1_FB2_BB1_IO_116,
    output wire        mb1_FA1_TB2_IO_115_mb1_FB2_BB1_IO_117,
    output wire        mb1_FA1_TB2_IO_116_mb1_FB2_BB1_IO_114,
    output wire        mb1_FA1_TB2_IO_117_mb1_FB2_BB1_IO_115,
    output wire        mb1_FA1_TB2_IO_118_mb1_FB2_BB1_IO_132,
    output wire        mb1_FA1_TB2_IO_119_mb1_FB2_BB1_IO_133,
    output wire        mb1_FA1_TB2_IO_120_mb1_FB2_BB1_IO_130,
    output wire        mb1_FA1_TB2_IO_121_mb1_FB2_BB1_IO_131,
    output wire        mb1_FA1_TB2_IO_122_mb1_FB2_BB1_IO_108,
    output wire        mb1_FA1_TB2_IO_123_mb1_FB2_BB1_IO_109,
    output wire        mb1_FA1_TB2_IO_124_mb1_FB2_BB1_IO_126,
    output wire        mb1_FA1_TB2_IO_125_mb1_FB2_BB1_IO_127,
    output wire        mb1_FA1_TB2_IO_126_mb1_FB2_BB1_IO_124,
    output wire        mb1_FA1_TB2_IO_127_mb1_FB2_BB1_IO_125,
    output wire        mb1_FA1_TB2_IO_130_mb1_FB2_BB1_IO_120,
    output wire        mb1_FA1_TB2_IO_131_mb1_FB2_BB1_IO_121,
    output wire        mb1_FA1_TB2_IO_132_mb1_FB2_BB1_IO_118,
    output wire        mb1_FA1_TB2_IO_133_mb1_FB2_BB1_IO_119,
    output wire        mb1_FA1_TB2_IO_134_mb1_FB2_BB1_IO_136,
    output wire        mb1_FA1_TB2_IO_136_mb1_FB2_BB1_IO_134,
    output wire        mb1_FA1_BA0_CLKIO_N_0_mb1_FB1_BA2_CLKIO_N_7,
    output wire        mb1_FA1_BA0_CLKIO_N_1_mb1_FB1_BA2_CLKIO_N_6,
    output wire        mb1_FA1_BA0_CLKIO_N_2_mb1_FB1_BA2_CLKIO_N_4,
    output wire        mb1_FA1_BA0_CLKIO_N_3_mb1_FB1_BA2_CLKIO_N_3,
    output wire        mb1_FA1_BA0_CLKIO_N_4_mb1_FB1_BA2_CLKIO_N_2,
    output wire        mb1_FA1_BA0_CLKIO_N_5_mb1_FB1_BA2_IO_010,
    output wire        mb1_FA1_BA0_CLKIO_N_6_mb1_FB1_BA2_CLKIO_N_1,
    output wire        mb1_FA1_BA0_CLKIO_N_7_mb1_FB1_BA2_CLKIO_N_0,
    output wire        mb1_FA1_BA0_CLKIO_P_0_mb1_FB1_BA2_CLKIO_P_7,
    output wire        mb1_FA1_BA0_CLKIO_P_1_mb1_FB1_BA2_CLKIO_P_6,
    output wire        mb1_FA1_BA0_CLKIO_P_2_mb1_FB1_BA2_CLKIO_P_4,
    output wire        mb1_FA1_BA0_CLKIO_P_3_mb1_FB1_BA2_CLKIO_P_3,
    output wire        mb1_FA1_BA0_CLKIO_P_4_mb1_FB1_BA2_CLKIO_P_2,
    output wire        mb1_FA1_BA0_CLKIO_P_5_mb1_FB1_BA2_IO_011,
    output wire        mb1_FA1_BA0_CLKIO_P_6_mb1_FB1_BA2_CLKIO_P_1,
    output wire        mb1_FA1_BA0_CLKIO_P_7_mb1_FB1_BA2_CLKIO_P_0,
    output wire        mb1_FA1_BA0_IO_004_mb1_FB1_BA2_IO_006,
    output wire        mb1_FA1_BA0_IO_005_mb1_FB1_BA2_IO_007,
    output wire        mb1_FA1_BA0_IO_006_mb1_FB1_BA2_IO_004,
    output wire        mb1_FA1_BA0_IO_007_mb1_FB1_BA2_IO_005,
    output wire        mb1_FA1_BA0_IO_008_mb1_FB1_BA2_IO_022,
    output wire        mb1_FA1_BA0_IO_009_mb1_FB1_BA2_IO_023,
    output wire        mb1_FA1_BA0_IO_010_mb1_FB1_BA2_CLKIO_N_5,
    output wire        mb1_FA1_BA0_IO_011_mb1_FB1_BA2_CLKIO_P_5,
    output wire        mb1_FA1_BA0_IO_012_mb1_FB1_BA2_IO_012,
    output wire        mb1_FA1_BA0_IO_013_mb1_FB1_BA2_IO_013,
    output wire        mb1_FA1_BA0_IO_014_mb1_FB1_BA2_IO_016,
    output wire        mb1_FA1_BA0_IO_015_mb1_FB1_BA2_IO_017,
    output wire        mb1_FA1_BA0_IO_016_mb1_FB1_BA2_IO_014,
    output wire        mb1_FA1_BA0_IO_017_mb1_FB1_BA2_IO_015,
    output wire        mb1_FA1_BA0_IO_018_mb1_FB1_BA2_IO_032,
    output wire        mb1_FA1_BA0_IO_019_mb1_FB1_BA2_IO_033,
    output wire        mb1_FA1_BA0_IO_020_mb1_FB1_BA2_IO_030,
    output wire        mb1_FA1_BA0_IO_021_mb1_FB1_BA2_IO_031,
    output wire        mb1_FA1_BA0_IO_022_mb1_FB1_BA2_IO_008,
    output wire        mb1_FA1_BA0_IO_023_mb1_FB1_BA2_IO_009,
    output wire        mb1_FA1_BA0_IO_024_mb1_FB1_BA2_IO_026,
    output wire        mb1_FA1_BA0_IO_025_mb1_FB1_BA2_IO_027,
    output wire        mb1_FA1_BA0_IO_026_mb1_FB1_BA2_IO_024,
    output wire        mb1_FA1_BA0_IO_027_mb1_FB1_BA2_IO_025,
    output wire        mb1_FA1_BA0_IO_028_mb1_FB1_BA2_IO_042,
    output wire        mb1_FA1_BA0_IO_029_mb1_FB1_BA2_IO_043,
    output wire        mb1_FA1_BA0_IO_030_mb1_FB1_BA2_IO_020,
    output wire        mb1_FA1_BA0_IO_031_mb1_FB1_BA2_IO_021,
    output wire        mb1_FA1_BA0_IO_032_mb1_FB1_BA2_IO_018,
    output wire        mb1_FA1_BA0_IO_033_mb1_FB1_BA2_IO_019,
    output wire        mb1_FA1_BA0_IO_034_mb1_FB1_BA2_IO_036,
    output wire        mb1_FA1_BA0_IO_035_mb1_FB1_BA2_IO_037,
    output wire        mb1_FA1_BA0_IO_036_mb1_FB1_BA2_IO_034,
    output wire        mb1_FA1_BA0_IO_037_mb1_FB1_BA2_IO_035,
    output wire        mb1_FA1_BA0_IO_038_mb1_FB1_BA2_IO_052,
    output wire        mb1_FA1_BA0_IO_039_mb1_FB1_BA2_IO_053,
    output wire        mb1_FA1_BA0_IO_040_mb1_FB1_BA2_IO_050,
    output wire        mb1_FA1_BA0_IO_041_mb1_FB1_BA2_IO_051,
    output wire        mb1_FA1_BA0_IO_042_mb1_FB1_BA2_IO_028,
    output wire        mb1_FA1_BA0_IO_043_mb1_FB1_BA2_IO_029,
    output wire        mb1_FA1_BA0_IO_044_mb1_FB1_BA2_IO_046,
    output wire        mb1_FA1_BA0_IO_045_mb1_FB1_BA2_IO_047,
    output wire        mb1_FA1_BA0_IO_046_mb1_FB1_BA2_IO_044,
    output wire        mb1_FA1_BA0_IO_047_mb1_FB1_BA2_IO_045,
    output wire        mb1_FA1_BA0_IO_048_mb1_FB1_BA2_IO_062,
    output wire        mb1_FA1_BA0_IO_049_mb1_FB1_BA2_IO_063,
    output wire        mb1_FA1_BA0_IO_050_mb1_FB1_BA2_IO_040,
    output wire        mb1_FA1_BA0_IO_051_mb1_FB1_BA2_IO_041,
    output wire        mb1_FA1_BA0_IO_052_mb1_FB1_BA2_IO_038,
    output wire        mb1_FA1_BA0_IO_053_mb1_FB1_BA2_IO_039,
    output wire        mb1_FA1_BA0_IO_054_mb1_FB1_BA2_IO_056,
    output wire        mb1_FA1_BA0_IO_055_mb1_FB1_BA2_IO_057,
    output wire        mb1_FA1_BA0_IO_056_mb1_FB1_BA2_IO_054,
    output wire        mb1_FA1_BA0_IO_057_mb1_FB1_BA2_IO_055,
    output wire        mb1_FA1_BA0_IO_058_mb1_FB1_BA2_IO_072,
    output wire        mb1_FA1_BA0_IO_059_mb1_FB1_BA2_IO_073,
    output wire        mb1_FA1_BA0_IO_060_mb1_FB1_BA2_IO_070,
    output wire        mb1_FA1_BA0_IO_061_mb1_FB1_BA2_IO_071,
    output wire        mb1_FA1_BA0_IO_062_mb1_FB1_BA2_IO_048,
    output wire        mb1_FA1_BA0_IO_063_mb1_FB1_BA2_IO_049,
    output wire        mb1_FA1_BA0_IO_064_mb1_FB1_BA2_IO_066,
    output wire        mb1_FA1_BA0_IO_065_mb1_FB1_BA2_IO_067,
    output wire        mb1_FA1_BA0_IO_066_mb1_FB1_BA2_IO_064,
    output wire        mb1_FA1_BA0_IO_067_mb1_FB1_BA2_IO_065,
    output wire        mb1_FA1_BA0_IO_068_mb1_FB1_BA2_IO_082,
    output wire        mb1_FA1_BA0_IO_069_mb1_FB1_BA2_IO_083,
    output wire        mb1_FA1_BA0_IO_070_mb1_FB1_BA2_IO_060,
    output wire        mb1_FA1_BA0_IO_071_mb1_FB1_BA2_IO_061,
    output wire        mb1_FA1_BA0_IO_072_mb1_FB1_BA2_IO_058,
    output wire        mb1_FA1_BA0_IO_073_mb1_FB1_BA2_IO_059,
    output wire        mb1_FA1_BA0_IO_074_mb1_FB1_BA2_IO_076,
    output wire        mb1_FA1_BA0_IO_075_mb1_FB1_BA2_IO_077,
    output wire        mb1_FA1_BA0_IO_076_mb1_FB1_BA2_IO_074,
    output wire        mb1_FA1_BA0_IO_077_mb1_FB1_BA2_IO_075,
    output wire        mb1_FA1_BA0_IO_078_mb1_FB1_BA2_IO_092,
    output wire        mb1_FA1_BA0_IO_079_mb1_FB1_BA2_IO_093,
    output wire        mb1_FA1_BA0_IO_080_mb1_FB1_BA2_IO_090,
    output wire        mb1_FA1_BA0_IO_081_mb1_FB1_BA2_IO_091,
    output wire        mb1_FA1_BA0_IO_082_mb1_FB1_BA2_IO_068,
    output wire        mb1_FA1_BA0_IO_083_mb1_FB1_BA2_IO_069,
    output wire        mb1_FA1_BA0_IO_084_mb1_FB1_BA2_IO_086,
    output wire        mb1_FA1_BA0_IO_085_mb1_FB1_BA2_IO_087,
    output wire        mb1_FA1_BA0_IO_086_mb1_FB1_BA2_IO_084,
    output wire        mb1_FA1_BA0_IO_087_mb1_FB1_BA2_IO_085,
    output wire        mb1_FA1_BA0_IO_088_mb1_FB1_BA2_IO_102,
    output wire        mb1_FA1_BA0_IO_089_mb1_FB1_BA2_IO_103,
    output wire        mb1_FA1_BA0_IO_090_mb1_FB1_BA2_IO_080,
    output wire        mb1_FA1_BA0_IO_091_mb1_FB1_BA2_IO_081,
    output wire        mb1_FA1_BA0_IO_092_mb1_FB1_BA2_IO_078,
    output wire        mb1_FA1_BA0_IO_093_mb1_FB1_BA2_IO_079,
    output wire        mb1_FA1_BA0_IO_094_mb1_FB1_BA2_IO_096,
    output wire        mb1_FA1_BA0_IO_095_mb1_FB1_BA2_IO_097,
    output wire        mb1_FA1_BA0_IO_096_mb1_FB1_BA2_IO_094,
    output wire        mb1_FA1_BA0_IO_097_mb1_FB1_BA2_IO_095,
    output wire        mb1_FA1_BA0_IO_098_mb1_FB1_BA2_IO_112,
    output wire        mb1_FA1_BA0_IO_099_mb1_FB1_BA2_IO_113,
    output wire        mb1_FA1_BA0_IO_100_mb1_FB1_BA2_IO_110,
    output wire        mb1_FA1_BA0_IO_101_mb1_FB1_BA2_IO_111,
    output wire        mb1_FA1_BA0_IO_102_mb1_FB1_BA2_IO_088,
    output wire        mb1_FA1_BA0_IO_103_mb1_FB1_BA2_IO_089,
    output wire        mb1_FA1_BA0_IO_104_mb1_FB1_BA2_IO_106,
    output wire        mb1_FA1_BA0_IO_105_mb1_FB1_BA2_IO_107,
    output wire        mb1_FA1_BA0_IO_106_mb1_FB1_BA2_IO_104,
    output wire        mb1_FA1_BA0_IO_107_mb1_FB1_BA2_IO_105,
    output wire        mb1_FA1_BA0_IO_108_mb1_FB1_BA2_IO_122,
    output wire        mb1_FA1_BA0_IO_109_mb1_FB1_BA2_IO_123,
    output wire        mb1_FA1_BA0_IO_110_mb1_FB1_BA2_IO_100,
    output wire        mb1_FA1_BA0_IO_111_mb1_FB1_BA2_IO_101,
    output wire        mb1_FA1_BA0_IO_112_mb1_FB1_BA2_IO_098,
    output wire        mb1_FA1_BA0_IO_113_mb1_FB1_BA2_IO_099,
    output wire        mb1_FA1_BA0_IO_114_mb1_FB1_BA2_IO_116,
    output wire        mb1_FA1_BA0_IO_115_mb1_FB1_BA2_IO_117,
    output wire        mb1_FA1_BA0_IO_116_mb1_FB1_BA2_IO_114,
    output wire        mb1_FA1_BA0_IO_117_mb1_FB1_BA2_IO_115,
    output wire        mb1_FA1_BA0_IO_118_mb1_FB1_BA2_IO_132,
    output wire        mb1_FA1_BA0_IO_119_mb1_FB1_BA2_IO_133,
    output wire        mb1_FA1_BA0_IO_120_mb1_FB1_BA2_IO_130,
    output wire        mb1_FA1_BA0_IO_121_mb1_FB1_BA2_IO_131,
    output wire        mb1_FA1_BA0_IO_122_mb1_FB1_BA2_IO_108,
    output wire        mb1_FA1_BA0_IO_123_mb1_FB1_BA2_IO_109,
    output wire        mb1_FA1_BA0_IO_124_mb1_FB1_BA2_IO_126,
    output wire        mb1_FA1_BA0_IO_125_mb1_FB1_BA2_IO_127,
    output wire        mb1_FA1_BA0_IO_126_mb1_FB1_BA2_IO_124,
    output wire        mb1_FA1_BA0_IO_127_mb1_FB1_BA2_IO_125,
    output wire        mb1_FA1_BA0_IO_130_mb1_FB1_BA2_IO_120,
    output wire        mb1_FA1_BA0_IO_131_mb1_FB1_BA2_IO_121,
    output wire        mb1_FA1_BA0_IO_132_mb1_FB1_BA2_IO_118,
    output wire        mb1_FA1_BA0_IO_133_mb1_FB1_BA2_IO_119,
    output wire        mb1_FA1_BA0_IO_134_mb1_FB1_BA2_IO_136,
    output wire        mb1_FA1_BA0_IO_136_mb1_FB1_BA2_IO_134,
    output wire        mb1_FA1_BA1_CLKIO_N_0_mb1_FA2_BB2_CLKIO_N_7,
    output wire        mb1_FA1_BA1_CLKIO_N_1_mb1_FA2_BB2_CLKIO_N_6,
    output wire        mb1_FA1_BA1_CLKIO_N_2_mb1_FA2_BB2_CLKIO_N_4,
    output wire        mb1_FA1_BA1_CLKIO_N_3_mb1_FA2_BB2_CLKIO_N_3,
    output wire        mb1_FA1_BA1_CLKIO_N_4_mb1_FA2_BB2_CLKIO_N_2,
    output wire        mb1_FA1_BA1_CLKIO_N_5_mb1_FA2_BB2_IO_010,
    output wire        mb1_FA1_BA1_CLKIO_N_6_mb1_FA2_BB2_CLKIO_N_1,
    output wire        mb1_FA1_BA1_CLKIO_N_7_mb1_FA2_BB2_CLKIO_N_0,
    output wire        mb1_FA1_BA1_CLKIO_P_0_mb1_FA2_BB2_CLKIO_P_7,
    output wire        mb1_FA1_BA1_CLKIO_P_1_mb1_FA2_BB2_CLKIO_P_6,
    output wire        mb1_FA1_BA1_CLKIO_P_2_mb1_FA2_BB2_CLKIO_P_4,
    output wire        mb1_FA1_BA1_CLKIO_P_3_mb1_FA2_BB2_CLKIO_P_3,
    output wire        mb1_FA1_BA1_CLKIO_P_4_mb1_FA2_BB2_CLKIO_P_2,
    output wire        mb1_FA1_BA1_CLKIO_P_5_mb1_FA2_BB2_IO_011,
    output wire        mb1_FA1_BA1_CLKIO_P_6_mb1_FA2_BB2_CLKIO_P_1,
    output wire        mb1_FA1_BA1_CLKIO_P_7_mb1_FA2_BB2_CLKIO_P_0,
    output wire        mb1_FA1_BA1_IO_004_mb1_FA2_BB2_IO_006,
    output wire        mb1_FA1_BA1_IO_005_mb1_FA2_BB2_IO_007,
    output wire        mb1_FA1_BA1_IO_006_mb1_FA2_BB2_IO_004,
    output wire        mb1_FA1_BA1_IO_007_mb1_FA2_BB2_IO_005,
    output wire        mb1_FA1_BA1_IO_008_mb1_FA2_BB2_IO_022,
    output wire        mb1_FA1_BA1_IO_009_mb1_FA2_BB2_IO_023,
    output wire        mb1_FA1_BA1_IO_010_mb1_FA2_BB2_CLKIO_N_5,
    output wire        mb1_FA1_BA1_IO_011_mb1_FA2_BB2_CLKIO_P_5,
    output wire        mb1_FA1_BA1_IO_012_mb1_FA2_BB2_IO_012,
    output wire        mb1_FA1_BA1_IO_013_mb1_FA2_BB2_IO_013,
    output wire        mb1_FA1_BA1_IO_014_mb1_FA2_BB2_IO_016,
    output wire        mb1_FA1_BA1_IO_015_mb1_FA2_BB2_IO_017,
    output wire        mb1_FA1_BA1_IO_016_mb1_FA2_BB2_IO_014,
    output wire        mb1_FA1_BA1_IO_017_mb1_FA2_BB2_IO_015,
    output wire        mb1_FA1_BA1_IO_018_mb1_FA2_BB2_IO_032,
    output wire        mb1_FA1_BA1_IO_019_mb1_FA2_BB2_IO_033,
    output wire        mb1_FA1_BA1_IO_020_mb1_FA2_BB2_IO_030,
    output wire        mb1_FA1_BA1_IO_021_mb1_FA2_BB2_IO_031,
    output wire        mb1_FA1_BA1_IO_022_mb1_FA2_BB2_IO_008,
    output wire        mb1_FA1_BA1_IO_023_mb1_FA2_BB2_IO_009,
    output wire        mb1_FA1_BA1_IO_024_mb1_FA2_BB2_IO_026,
    output wire        mb1_FA1_BA1_IO_025_mb1_FA2_BB2_IO_027,
    output wire        mb1_FA1_BA1_IO_026_mb1_FA2_BB2_IO_024,
    output wire        mb1_FA1_BA1_IO_027_mb1_FA2_BB2_IO_025,
    output wire        mb1_FA1_BA1_IO_028_mb1_FA2_BB2_IO_042,
    output wire        mb1_FA1_BA1_IO_029_mb1_FA2_BB2_IO_043,
    output wire        mb1_FA1_BA1_IO_030_mb1_FA2_BB2_IO_020,
    output wire        mb1_FA1_BA1_IO_031_mb1_FA2_BB2_IO_021,
    output wire        mb1_FA1_BA1_IO_032_mb1_FA2_BB2_IO_018,
    output wire        mb1_FA1_BA1_IO_033_mb1_FA2_BB2_IO_019,
    output wire        mb1_FA1_BA1_IO_034_mb1_FA2_BB2_IO_036,
    output wire        mb1_FA1_BA1_IO_035_mb1_FA2_BB2_IO_037,
    output wire        mb1_FA1_BA1_IO_036_mb1_FA2_BB2_IO_034,
    output wire        mb1_FA1_BA1_IO_037_mb1_FA2_BB2_IO_035,
    output wire        mb1_FA1_BA1_IO_038_mb1_FA2_BB2_IO_052,
    output wire        mb1_FA1_BA1_IO_039_mb1_FA2_BB2_IO_053,
    output wire        mb1_FA1_BA1_IO_040_mb1_FA2_BB2_IO_050,
    output wire        mb1_FA1_BA1_IO_041_mb1_FA2_BB2_IO_051,
    output wire        mb1_FA1_BA1_IO_042_mb1_FA2_BB2_IO_028,
    output wire        mb1_FA1_BA1_IO_043_mb1_FA2_BB2_IO_029,
    output wire        mb1_FA1_BA1_IO_044_mb1_FA2_BB2_IO_046,
    output wire        mb1_FA1_BA1_IO_045_mb1_FA2_BB2_IO_047,
    output wire        mb1_FA1_BA1_IO_046_mb1_FA2_BB2_IO_044,
    output wire        mb1_FA1_BA1_IO_047_mb1_FA2_BB2_IO_045,
    output wire        mb1_FA1_BA1_IO_048_mb1_FA2_BB2_IO_062,
    output wire        mb1_FA1_BA1_IO_049_mb1_FA2_BB2_IO_063,
    output wire        mb1_FA1_BA1_IO_050_mb1_FA2_BB2_IO_040,
    output wire        mb1_FA1_BA1_IO_051_mb1_FA2_BB2_IO_041,
    output wire        mb1_FA1_BA1_IO_052_mb1_FA2_BB2_IO_038,
    output wire        mb1_FA1_BA1_IO_053_mb1_FA2_BB2_IO_039,
    output wire        mb1_FA1_BA1_IO_054_mb1_FA2_BB2_IO_056,
    output wire        mb1_FA1_BA1_IO_055_mb1_FA2_BB2_IO_057,
    output wire        mb1_FA1_BA1_IO_056_mb1_FA2_BB2_IO_054,
    output wire        mb1_FA1_BA1_IO_057_mb1_FA2_BB2_IO_055,
    output wire        mb1_FA1_BA1_IO_058_mb1_FA2_BB2_IO_072,
    output wire        mb1_FA1_BA1_IO_059_mb1_FA2_BB2_IO_073,
    output wire        mb1_FA1_BA1_IO_060_mb1_FA2_BB2_IO_070,
    output wire        mb1_FA1_BA1_IO_061_mb1_FA2_BB2_IO_071,
    output wire        mb1_FA1_BA1_IO_062_mb1_FA2_BB2_IO_048,
    output wire        mb1_FA1_BA1_IO_063_mb1_FA2_BB2_IO_049,
    output wire        mb1_FA1_BA1_IO_064_mb1_FA2_BB2_IO_066,
    output wire        mb1_FA1_BA1_IO_065_mb1_FA2_BB2_IO_067,
    output wire        mb1_FA1_BA1_IO_066_mb1_FA2_BB2_IO_064,
    output wire        mb1_FA1_BA1_IO_067_mb1_FA2_BB2_IO_065,
    output wire        mb1_FA1_BA1_IO_068_mb1_FA2_BB2_IO_082,
    output wire        mb1_FA1_BA1_IO_069_mb1_FA2_BB2_IO_083,
    output wire        mb1_FA1_BA1_IO_070_mb1_FA2_BB2_IO_060,
    output wire        mb1_FA1_BA1_IO_071_mb1_FA2_BB2_IO_061,
    output wire        mb1_FA1_BA1_IO_072_mb1_FA2_BB2_IO_058,
    output wire        mb1_FA1_BA1_IO_073_mb1_FA2_BB2_IO_059,
    output wire        mb1_FA1_BA1_IO_074_mb1_FA2_BB2_IO_076,
    output wire        mb1_FA1_BA1_IO_075_mb1_FA2_BB2_IO_077,
    output wire        mb1_FA1_BA1_IO_076_mb1_FA2_BB2_IO_074,
    output wire        mb1_FA1_BA1_IO_077_mb1_FA2_BB2_IO_075,
    output wire        mb1_FA1_BA1_IO_078_mb1_FA2_BB2_IO_092,
    output wire        mb1_FA1_BA1_IO_079_mb1_FA2_BB2_IO_093,
    output wire        mb1_FA1_BA1_IO_080_mb1_FA2_BB2_IO_090,
    output wire        mb1_FA1_BA1_IO_081_mb1_FA2_BB2_IO_091,
    output wire        mb1_FA1_BA1_IO_082_mb1_FA2_BB2_IO_068,
    output wire        mb1_FA1_BA1_IO_083_mb1_FA2_BB2_IO_069,
    output wire        mb1_FA1_BA1_IO_084_mb1_FA2_BB2_IO_086,
    output wire        mb1_FA1_BA1_IO_085_mb1_FA2_BB2_IO_087,
    output wire        mb1_FA1_BA1_IO_086_mb1_FA2_BB2_IO_084,
    output wire        mb1_FA1_BA1_IO_087_mb1_FA2_BB2_IO_085,
    output wire        mb1_FA1_BA1_IO_088_mb1_FA2_BB2_IO_102,
    output wire        mb1_FA1_BA1_IO_089_mb1_FA2_BB2_IO_103,
    output wire        mb1_FA1_BA1_IO_090_mb1_FA2_BB2_IO_080,
    output wire        mb1_FA1_BA1_IO_091_mb1_FA2_BB2_IO_081,
    output wire        mb1_FA1_BA1_IO_092_mb1_FA2_BB2_IO_078,
    output wire        mb1_FA1_BA1_IO_093_mb1_FA2_BB2_IO_079,
    output wire        mb1_FA1_BA1_IO_094_mb1_FA2_BB2_IO_096,
    output wire        mb1_FA1_BA1_IO_095_mb1_FA2_BB2_IO_097,
    output wire        mb1_FA1_BA1_IO_096_mb1_FA2_BB2_IO_094,
    output wire        mb1_FA1_BA1_IO_097_mb1_FA2_BB2_IO_095,
    output wire        mb1_FA1_BA1_IO_098_mb1_FA2_BB2_IO_112,
    output wire        mb1_FA1_BA1_IO_099_mb1_FA2_BB2_IO_113,
    output wire        mb1_FA1_BA1_IO_100_mb1_FA2_BB2_IO_110,
    output wire        mb1_FA1_BA1_IO_101_mb1_FA2_BB2_IO_111,
    output wire        mb1_FA1_BA1_IO_102_mb1_FA2_BB2_IO_088,
    output wire        mb1_FA1_BA1_IO_103_mb1_FA2_BB2_IO_089,
    output wire        mb1_FA1_BA1_IO_104_mb1_FA2_BB2_IO_106,
    output wire        mb1_FA1_BA1_IO_105_mb1_FA2_BB2_IO_107,
    output wire        mb1_FA1_BA1_IO_106_mb1_FA2_BB2_IO_104,
    output wire        mb1_FA1_BA1_IO_107_mb1_FA2_BB2_IO_105,
    output wire        mb1_FA1_BA1_IO_108_mb1_FA2_BB2_IO_122,
    output wire        mb1_FA1_BA1_IO_109_mb1_FA2_BB2_IO_123,
    output wire        mb1_FA1_BA1_IO_110_mb1_FA2_BB2_IO_100,
    output wire        mb1_FA1_BA1_IO_111_mb1_FA2_BB2_IO_101,
    output wire        mb1_FA1_BA1_IO_112_mb1_FA2_BB2_IO_098,
    output wire        mb1_FA1_BA1_IO_113_mb1_FA2_BB2_IO_099,
    output wire        mb1_FA1_BA1_IO_114_mb1_FA2_BB2_IO_116,
    output wire        mb1_FA1_BA1_IO_115_mb1_FA2_BB2_IO_117,
    output wire        mb1_FA1_BA1_IO_116_mb1_FA2_BB2_IO_114,
    output wire        mb1_FA1_BA1_IO_117_mb1_FA2_BB2_IO_115,
    output wire        mb1_FA1_BA1_IO_118_mb1_FA2_BB2_IO_132,
    output wire        mb1_FA1_BA1_IO_119_mb1_FA2_BB2_IO_133,
    output wire        mb1_FA1_BA1_IO_120_mb1_FA2_BB2_IO_130,
    output wire        mb1_FA1_BA1_IO_121_mb1_FA2_BB2_IO_131,
    output wire        mb1_FA1_BA1_IO_122_mb1_FA2_BB2_IO_108,
    output wire        mb1_FA1_BA1_IO_123_mb1_FA2_BB2_IO_109,
    output wire        mb1_FA1_BA1_IO_124_mb1_FA2_BB2_IO_126,
    output wire        mb1_FA1_BA1_IO_125_mb1_FA2_BB2_IO_127,
    output wire        mb1_FA1_BA1_IO_126_mb1_FA2_BB2_IO_124,
    output wire        mb1_FA1_BA1_IO_127_mb1_FA2_BB2_IO_125,
    output wire        mb1_FA1_BA1_IO_130_mb1_FA2_BB2_IO_120,
    output wire        mb1_FA1_BA1_IO_131_mb1_FA2_BB2_IO_121,
    output wire        mb1_FA1_BA1_IO_132_mb1_FA2_BB2_IO_118,
    output wire        mb1_FA1_BA1_IO_133_mb1_FA2_BB2_IO_119,
    output wire        mb1_FA1_BA1_IO_134_mb1_FA2_BB2_IO_136,
    output wire        mb1_FA1_BA1_IO_136_mb1_FA2_BB2_IO_134,
    output wire        mb1_FA1_BA2_CLKIO_N_0_mb1_FB1_BB0_CLKIO_N_7,
    output wire        mb1_FA1_BA2_CLKIO_N_1_mb1_FB1_BB0_CLKIO_N_6,
    output wire        mb1_FA1_BA2_CLKIO_N_2_mb1_FB1_BB0_CLKIO_N_4,
    output wire        mb1_FA1_BA2_CLKIO_N_3_mb1_FB1_BB0_CLKIO_N_3,
    output wire        mb1_FA1_BA2_CLKIO_N_4_mb1_FB1_BB0_CLKIO_N_2,
    output wire        mb1_FA1_BA2_CLKIO_N_5_mb1_FB1_BB0_IO_010,
    output wire        mb1_FA1_BA2_CLKIO_N_6_mb1_FB1_BB0_CLKIO_N_1,
    output wire        mb1_FA1_BA2_CLKIO_N_7_mb1_FB1_BB0_CLKIO_N_0,
    output wire        mb1_FA1_BA2_CLKIO_P_0_mb1_FB1_BB0_CLKIO_P_7,
    output wire        mb1_FA1_BA2_CLKIO_P_1_mb1_FB1_BB0_CLKIO_P_6,
    output wire        mb1_FA1_BA2_CLKIO_P_2_mb1_FB1_BB0_CLKIO_P_4,
    output wire        mb1_FA1_BA2_CLKIO_P_3_mb1_FB1_BB0_CLKIO_P_3,
    output wire        mb1_FA1_BA2_CLKIO_P_4_mb1_FB1_BB0_CLKIO_P_2,
    output wire        mb1_FA1_BA2_CLKIO_P_5_mb1_FB1_BB0_IO_011,
    output wire        mb1_FA1_BA2_CLKIO_P_6_mb1_FB1_BB0_CLKIO_P_1,
    output wire        mb1_FA1_BA2_CLKIO_P_7_mb1_FB1_BB0_CLKIO_P_0,
    output wire        mb1_FA1_BA2_IO_004_mb1_FB1_BB0_IO_006,
    output wire        mb1_FA1_BA2_IO_005_mb1_FB1_BB0_IO_007,
    output wire        mb1_FA1_BA2_IO_006_mb1_FB1_BB0_IO_004,
    output wire        mb1_FA1_BA2_IO_007_mb1_FB1_BB0_IO_005,
    output wire        mb1_FA1_BA2_IO_008_mb1_FB1_BB0_IO_022,
    output wire        mb1_FA1_BA2_IO_009_mb1_FB1_BB0_IO_023,
    output wire        mb1_FA1_BA2_IO_010_mb1_FB1_BB0_CLKIO_N_5,
    output wire        mb1_FA1_BA2_IO_011_mb1_FB1_BB0_CLKIO_P_5,
    output wire        mb1_FA1_BA2_IO_012_mb1_FB1_BB0_IO_012,
    output wire        mb1_FA1_BA2_IO_013_mb1_FB1_BB0_IO_013,
    output wire        mb1_FA1_BA2_IO_014_mb1_FB1_BB0_IO_016,
    output wire        mb1_FA1_BA2_IO_015_mb1_FB1_BB0_IO_017,
    output wire        mb1_FA1_BA2_IO_016_mb1_FB1_BB0_IO_014,
    output wire        mb1_FA1_BA2_IO_017_mb1_FB1_BB0_IO_015,
    output wire        mb1_FA1_BA2_IO_018_mb1_FB1_BB0_IO_032,
    output wire        mb1_FA1_BA2_IO_019_mb1_FB1_BB0_IO_033,
    output wire        mb1_FA1_BA2_IO_020_mb1_FB1_BB0_IO_030,
    output wire        mb1_FA1_BA2_IO_021_mb1_FB1_BB0_IO_031,
    output wire        mb1_FA1_BA2_IO_022_mb1_FB1_BB0_IO_008,
    output wire        mb1_FA1_BA2_IO_023_mb1_FB1_BB0_IO_009,
    output wire        mb1_FA1_BA2_IO_024_mb1_FB1_BB0_IO_026,
    output wire        mb1_FA1_BA2_IO_025_mb1_FB1_BB0_IO_027,
    output wire        mb1_FA1_BA2_IO_026_mb1_FB1_BB0_IO_024,
    output wire        mb1_FA1_BA2_IO_027_mb1_FB1_BB0_IO_025,
    output wire        mb1_FA1_BA2_IO_028_mb1_FB1_BB0_IO_042,
    output wire        mb1_FA1_BA2_IO_029_mb1_FB1_BB0_IO_043,
    output wire        mb1_FA1_BA2_IO_030_mb1_FB1_BB0_IO_020,
    output wire        mb1_FA1_BA2_IO_031_mb1_FB1_BB0_IO_021,
    output wire        mb1_FA1_BA2_IO_032_mb1_FB1_BB0_IO_018,
    output wire        mb1_FA1_BA2_IO_033_mb1_FB1_BB0_IO_019,
    output wire        mb1_FA1_BA2_IO_034_mb1_FB1_BB0_IO_036,
    output wire        mb1_FA1_BA2_IO_035_mb1_FB1_BB0_IO_037,
    output wire        mb1_FA1_BA2_IO_036_mb1_FB1_BB0_IO_034,
    output wire        mb1_FA1_BA2_IO_037_mb1_FB1_BB0_IO_035,
    output wire        mb1_FA1_BA2_IO_038_mb1_FB1_BB0_IO_052,
    output wire        mb1_FA1_BA2_IO_039_mb1_FB1_BB0_IO_053,
    output wire        mb1_FA1_BA2_IO_040_mb1_FB1_BB0_IO_050,
    output wire        mb1_FA1_BA2_IO_041_mb1_FB1_BB0_IO_051,
    output wire        mb1_FA1_BA2_IO_042_mb1_FB1_BB0_IO_028,
    output wire        mb1_FA1_BA2_IO_043_mb1_FB1_BB0_IO_029,
    output wire        mb1_FA1_BA2_IO_044_mb1_FB1_BB0_IO_046,
    output wire        mb1_FA1_BA2_IO_045_mb1_FB1_BB0_IO_047,
    output wire        mb1_FA1_BA2_IO_046_mb1_FB1_BB0_IO_044,
    output wire        mb1_FA1_BA2_IO_047_mb1_FB1_BB0_IO_045,
    output wire        mb1_FA1_BA2_IO_048_mb1_FB1_BB0_IO_062,
    output wire        mb1_FA1_BA2_IO_049_mb1_FB1_BB0_IO_063,
    output wire        mb1_FA1_BA2_IO_050_mb1_FB1_BB0_IO_040,
    output wire        mb1_FA1_BA2_IO_051_mb1_FB1_BB0_IO_041,
    output wire        mb1_FA1_BA2_IO_052_mb1_FB1_BB0_IO_038,
    output wire        mb1_FA1_BA2_IO_053_mb1_FB1_BB0_IO_039,
    output wire        mb1_FA1_BA2_IO_054_mb1_FB1_BB0_IO_056,
    output wire        mb1_FA1_BA2_IO_055_mb1_FB1_BB0_IO_057,
    output wire        mb1_FA1_BA2_IO_056_mb1_FB1_BB0_IO_054,
    output wire        mb1_FA1_BA2_IO_057_mb1_FB1_BB0_IO_055,
    output wire        mb1_FA1_BA2_IO_058_mb1_FB1_BB0_IO_072,
    output wire        mb1_FA1_BA2_IO_059_mb1_FB1_BB0_IO_073,
    output wire        mb1_FA1_BA2_IO_060_mb1_FB1_BB0_IO_070,
    output wire        mb1_FA1_BA2_IO_061_mb1_FB1_BB0_IO_071,
    output wire        mb1_FA1_BA2_IO_062_mb1_FB1_BB0_IO_048,
    output wire        mb1_FA1_BA2_IO_063_mb1_FB1_BB0_IO_049,
    output wire        mb1_FA1_BA2_IO_064_mb1_FB1_BB0_IO_066,
    output wire        mb1_FA1_BA2_IO_065_mb1_FB1_BB0_IO_067,
    output wire        mb1_FA1_BA2_IO_066_mb1_FB1_BB0_IO_064,
    output wire        mb1_FA1_BA2_IO_067_mb1_FB1_BB0_IO_065,
    output wire        mb1_FA1_BA2_IO_068_mb1_FB1_BB0_IO_082,
    output wire        mb1_FA1_BA2_IO_069_mb1_FB1_BB0_IO_083,
    output wire        mb1_FA1_BA2_IO_070_mb1_FB1_BB0_IO_060,
    output wire        mb1_FA1_BA2_IO_071_mb1_FB1_BB0_IO_061,
    output wire        mb1_FA1_BA2_IO_072_mb1_FB1_BB0_IO_058,
    output wire        mb1_FA1_BA2_IO_073_mb1_FB1_BB0_IO_059,
    output wire        mb1_FA1_BA2_IO_074_mb1_FB1_BB0_IO_076,
    output wire        mb1_FA1_BA2_IO_075_mb1_FB1_BB0_IO_077,
    output wire        mb1_FA1_BA2_IO_076_mb1_FB1_BB0_IO_074,
    output wire        mb1_FA1_BA2_IO_077_mb1_FB1_BB0_IO_075,
    output wire        mb1_FA1_BA2_IO_078_mb1_FB1_BB0_IO_092,
    output wire        mb1_FA1_BA2_IO_079_mb1_FB1_BB0_IO_093,
    output wire        mb1_FA1_BA2_IO_080_mb1_FB1_BB0_IO_090,
    output wire        mb1_FA1_BA2_IO_081_mb1_FB1_BB0_IO_091,
    output wire        mb1_FA1_BA2_IO_082_mb1_FB1_BB0_IO_068,
    output wire        mb1_FA1_BA2_IO_083_mb1_FB1_BB0_IO_069,
    output wire        mb1_FA1_BA2_IO_084_mb1_FB1_BB0_IO_086,
    output wire        mb1_FA1_BA2_IO_085_mb1_FB1_BB0_IO_087,
    output wire        mb1_FA1_BA2_IO_086_mb1_FB1_BB0_IO_084,
    output wire        mb1_FA1_BA2_IO_087_mb1_FB1_BB0_IO_085,
    output wire        mb1_FA1_BA2_IO_088_mb1_FB1_BB0_IO_102,
    output wire        mb1_FA1_BA2_IO_089_mb1_FB1_BB0_IO_103,
    output wire        mb1_FA1_BA2_IO_090_mb1_FB1_BB0_IO_080,
    output wire        mb1_FA1_BA2_IO_091_mb1_FB1_BB0_IO_081,
    output wire        mb1_FA1_BA2_IO_092_mb1_FB1_BB0_IO_078,
    output wire        mb1_FA1_BA2_IO_093_mb1_FB1_BB0_IO_079,
    output wire        mb1_FA1_BA2_IO_094_mb1_FB1_BB0_IO_096,
    output wire        mb1_FA1_BA2_IO_095_mb1_FB1_BB0_IO_097,
    output wire        mb1_FA1_BA2_IO_096_mb1_FB1_BB0_IO_094,
    output wire        mb1_FA1_BA2_IO_097_mb1_FB1_BB0_IO_095,
    output wire        mb1_FA1_BA2_IO_098_mb1_FB1_BB0_IO_112,
    output wire        mb1_FA1_BA2_IO_099_mb1_FB1_BB0_IO_113,
    output wire        mb1_FA1_BA2_IO_100_mb1_FB1_BB0_IO_110,
    output wire        mb1_FA1_BA2_IO_101_mb1_FB1_BB0_IO_111,
    output wire        mb1_FA1_BA2_IO_102_mb1_FB1_BB0_IO_088,
    output wire        mb1_FA1_BA2_IO_103_mb1_FB1_BB0_IO_089,
    output wire        mb1_FA1_BA2_IO_104_mb1_FB1_BB0_IO_106,
    output wire        mb1_FA1_BA2_IO_105_mb1_FB1_BB0_IO_107,
    output wire        mb1_FA1_BA2_IO_106_mb1_FB1_BB0_IO_104,
    output wire        mb1_FA1_BA2_IO_107_mb1_FB1_BB0_IO_105,
    output wire        mb1_FA1_BA2_IO_108_mb1_FB1_BB0_IO_122,
    output wire        mb1_FA1_BA2_IO_109_mb1_FB1_BB0_IO_123,
    output wire        mb1_FA1_BA2_IO_110_mb1_FB1_BB0_IO_100,
    output wire        mb1_FA1_BA2_IO_111_mb1_FB1_BB0_IO_101,
    output wire        mb1_FA1_BA2_IO_112_mb1_FB1_BB0_IO_098,
    output wire        mb1_FA1_BA2_IO_113_mb1_FB1_BB0_IO_099,
    output wire        mb1_FA1_BA2_IO_114_mb1_FB1_BB0_IO_116,
    output wire        mb1_FA1_BA2_IO_115_mb1_FB1_BB0_IO_117,
    output wire        mb1_FA1_BA2_IO_116_mb1_FB1_BB0_IO_114,
    output wire        mb1_FA1_BA2_IO_117_mb1_FB1_BB0_IO_115,
    output wire        mb1_FA1_BA2_IO_118_mb1_FB1_BB0_IO_132,
    output wire        mb1_FA1_BA2_IO_119_mb1_FB1_BB0_IO_133,
    output wire        mb1_FA1_BA2_IO_120_mb1_FB1_BB0_IO_130,
    output wire        mb1_FA1_BA2_IO_121_mb1_FB1_BB0_IO_131,
    output wire        mb1_FA1_BA2_IO_122_mb1_FB1_BB0_IO_108,
    output wire        mb1_FA1_BA2_IO_123_mb1_FB1_BB0_IO_109,
    output wire        mb1_FA1_BA2_IO_124_mb1_FB1_BB0_IO_126,
    output wire        mb1_FA1_BA2_IO_125_mb1_FB1_BB0_IO_127,
    output wire        mb1_FA1_BA2_IO_126_mb1_FB1_BB0_IO_124,
    output wire        mb1_FA1_BA2_IO_127_mb1_FB1_BB0_IO_125,
    output wire        mb1_FA1_BA2_IO_130_mb1_FB1_BB0_IO_120,
    output wire        mb1_FA1_BA2_IO_131_mb1_FB1_BB0_IO_121,
    output wire        mb1_FA1_BA2_IO_132_mb1_FB1_BB0_IO_118,
    output wire        mb1_FA1_BA2_IO_133_mb1_FB1_BB0_IO_119,
    output wire        mb1_FA1_BA2_IO_134_mb1_FB1_BB0_IO_136,
    output wire        mb1_FA1_BA2_IO_136_mb1_FB1_BB0_IO_134,
    output wire        mb1_FA1_BB0_CLKIO_N_0_mb1_FB1_BB2_CLKIO_N_7,
    output wire        mb1_FA1_BB0_CLKIO_N_1_mb1_FB1_BB2_CLKIO_N_6,
    output wire        mb1_FA1_BB0_CLKIO_N_2_mb1_FB1_BB2_CLKIO_N_4,
    output wire        mb1_FA1_BB0_CLKIO_N_3_mb1_FB1_BB2_CLKIO_N_3,
    output wire        mb1_FA1_BB0_CLKIO_N_4_mb1_FB1_BB2_CLKIO_N_2,
    output wire        mb1_FA1_BB0_CLKIO_N_5_mb1_FB1_BB2_IO_010,
    output wire        mb1_FA1_BB0_CLKIO_N_6_mb1_FB1_BB2_CLKIO_N_1,
    output wire        mb1_FA1_BB0_CLKIO_N_7_mb1_FB1_BB2_CLKIO_N_0,
    output wire        mb1_FA1_BB0_CLKIO_P_0_mb1_FB1_BB2_CLKIO_P_7,
    output wire        mb1_FA1_BB0_CLKIO_P_1_mb1_FB1_BB2_CLKIO_P_6,
    output wire        mb1_FA1_BB0_CLKIO_P_2_mb1_FB1_BB2_CLKIO_P_4,
    output wire        mb1_FA1_BB0_CLKIO_P_3_mb1_FB1_BB2_CLKIO_P_3,
    output wire        mb1_FA1_BB0_CLKIO_P_4_mb1_FB1_BB2_CLKIO_P_2,
    output wire        mb1_FA1_BB0_CLKIO_P_5_mb1_FB1_BB2_IO_011,
    output wire        mb1_FA1_BB0_CLKIO_P_6_mb1_FB1_BB2_CLKIO_P_1,
    output wire        mb1_FA1_BB0_CLKIO_P_7_mb1_FB1_BB2_CLKIO_P_0,
    output wire        mb1_FA1_BB0_IO_004_mb1_FB1_BB2_IO_006,
    output wire        mb1_FA1_BB0_IO_005_mb1_FB1_BB2_IO_007,
    output wire        mb1_FA1_BB0_IO_006_mb1_FB1_BB2_IO_004,
    output wire        mb1_FA1_BB0_IO_007_mb1_FB1_BB2_IO_005,
    output wire        mb1_FA1_BB0_IO_008_mb1_FB1_BB2_IO_022,
    output wire        mb1_FA1_BB0_IO_009_mb1_FB1_BB2_IO_023,
    output wire        mb1_FA1_BB0_IO_010_mb1_FB1_BB2_CLKIO_N_5,
    output wire        mb1_FA1_BB0_IO_011_mb1_FB1_BB2_CLKIO_P_5,
    output wire        mb1_FA1_BB0_IO_012_mb1_FB1_BB2_IO_012,
    output wire        mb1_FA1_BB0_IO_013_mb1_FB1_BB2_IO_013,
    output wire        mb1_FA1_BB0_IO_014_mb1_FB1_BB2_IO_016,
    output wire        mb1_FA1_BB0_IO_015_mb1_FB1_BB2_IO_017,
    output wire        mb1_FA1_BB0_IO_016_mb1_FB1_BB2_IO_014,
    output wire        mb1_FA1_BB0_IO_017_mb1_FB1_BB2_IO_015,
    output wire        mb1_FA1_BB0_IO_018_mb1_FB1_BB2_IO_032,
    output wire        mb1_FA1_BB0_IO_019_mb1_FB1_BB2_IO_033,
    output wire        mb1_FA1_BB0_IO_020_mb1_FB1_BB2_IO_030,
    output wire        mb1_FA1_BB0_IO_021_mb1_FB1_BB2_IO_031,
    output wire        mb1_FA1_BB0_IO_022_mb1_FB1_BB2_IO_008,
    output wire        mb1_FA1_BB0_IO_023_mb1_FB1_BB2_IO_009,
    output wire        mb1_FA1_BB0_IO_024_mb1_FB1_BB2_IO_026,
    output wire        mb1_FA1_BB0_IO_025_mb1_FB1_BB2_IO_027,
    output wire        mb1_FA1_BB0_IO_026_mb1_FB1_BB2_IO_024,
    output wire        mb1_FA1_BB0_IO_027_mb1_FB1_BB2_IO_025,
    output wire        mb1_FA1_BB0_IO_028_mb1_FB1_BB2_IO_042,
    output wire        mb1_FA1_BB0_IO_029_mb1_FB1_BB2_IO_043,
    output wire        mb1_FA1_BB0_IO_030_mb1_FB1_BB2_IO_020,
    output wire        mb1_FA1_BB0_IO_031_mb1_FB1_BB2_IO_021,
    output wire        mb1_FA1_BB0_IO_032_mb1_FB1_BB2_IO_018,
    output wire        mb1_FA1_BB0_IO_033_mb1_FB1_BB2_IO_019,
    output wire        mb1_FA1_BB0_IO_034_mb1_FB1_BB2_IO_036,
    output wire        mb1_FA1_BB0_IO_035_mb1_FB1_BB2_IO_037,
    output wire        mb1_FA1_BB0_IO_036_mb1_FB1_BB2_IO_034,
    output wire        mb1_FA1_BB0_IO_037_mb1_FB1_BB2_IO_035,
    output wire        mb1_FA1_BB0_IO_038_mb1_FB1_BB2_IO_052,
    output wire        mb1_FA1_BB0_IO_039_mb1_FB1_BB2_IO_053,
    output wire        mb1_FA1_BB0_IO_040_mb1_FB1_BB2_IO_050,
    output wire        mb1_FA1_BB0_IO_041_mb1_FB1_BB2_IO_051,
    output wire        mb1_FA1_BB0_IO_042_mb1_FB1_BB2_IO_028,
    output wire        mb1_FA1_BB0_IO_043_mb1_FB1_BB2_IO_029,
    output wire        mb1_FA1_BB0_IO_044_mb1_FB1_BB2_IO_046,
    output wire        mb1_FA1_BB0_IO_045_mb1_FB1_BB2_IO_047,
    output wire        mb1_FA1_BB0_IO_046_mb1_FB1_BB2_IO_044,
    output wire        mb1_FA1_BB0_IO_047_mb1_FB1_BB2_IO_045,
    output wire        mb1_FA1_BB0_IO_048_mb1_FB1_BB2_IO_062,
    output wire        mb1_FA1_BB0_IO_049_mb1_FB1_BB2_IO_063,
    output wire        mb1_FA1_BB0_IO_050_mb1_FB1_BB2_IO_040,
    output wire        mb1_FA1_BB0_IO_051_mb1_FB1_BB2_IO_041,
    output wire        mb1_FA1_BB0_IO_052_mb1_FB1_BB2_IO_038,
    output wire        mb1_FA1_BB0_IO_053_mb1_FB1_BB2_IO_039,
    output wire        mb1_FA1_BB0_IO_054_mb1_FB1_BB2_IO_056,
    output wire        mb1_FA1_BB0_IO_055_mb1_FB1_BB2_IO_057,
    output wire        mb1_FA1_BB0_IO_056_mb1_FB1_BB2_IO_054,
    output wire        mb1_FA1_BB0_IO_057_mb1_FB1_BB2_IO_055,
    output wire        mb1_FA1_BB0_IO_058_mb1_FB1_BB2_IO_072,
    output wire        mb1_FA1_BB0_IO_059_mb1_FB1_BB2_IO_073,
    output wire        mb1_FA1_BB0_IO_060_mb1_FB1_BB2_IO_070,
    output wire        mb1_FA1_BB0_IO_061_mb1_FB1_BB2_IO_071,
    output wire        mb1_FA1_BB0_IO_062_mb1_FB1_BB2_IO_048,
    output wire        mb1_FA1_BB0_IO_063_mb1_FB1_BB2_IO_049,
    output wire        mb1_FA1_BB0_IO_064_mb1_FB1_BB2_IO_066,
    output wire        mb1_FA1_BB0_IO_065_mb1_FB1_BB2_IO_067,
    output wire        mb1_FA1_BB0_IO_066_mb1_FB1_BB2_IO_064,
    output wire        mb1_FA1_BB0_IO_067_mb1_FB1_BB2_IO_065,
    output wire        mb1_FA1_BB0_IO_068_mb1_FB1_BB2_IO_082,
    output wire        mb1_FA1_BB0_IO_069_mb1_FB1_BB2_IO_083,
    output wire        mb1_FA1_BB0_IO_070_mb1_FB1_BB2_IO_060,
    output wire        mb1_FA1_BB0_IO_071_mb1_FB1_BB2_IO_061,
    output wire        mb1_FA1_BB0_IO_072_mb1_FB1_BB2_IO_058,
    output wire        mb1_FA1_BB0_IO_073_mb1_FB1_BB2_IO_059,
    output wire        mb1_FA1_BB0_IO_074_mb1_FB1_BB2_IO_076,
    output wire        mb1_FA1_BB0_IO_075_mb1_FB1_BB2_IO_077,
    output wire        mb1_FA1_BB0_IO_076_mb1_FB1_BB2_IO_074,
    output wire        mb1_FA1_BB0_IO_077_mb1_FB1_BB2_IO_075,
    output wire        mb1_FA1_BB0_IO_078_mb1_FB1_BB2_IO_092,
    output wire        mb1_FA1_BB0_IO_079_mb1_FB1_BB2_IO_093,
    output wire        mb1_FA1_BB0_IO_080_mb1_FB1_BB2_IO_090,
    output wire        mb1_FA1_BB0_IO_081_mb1_FB1_BB2_IO_091,
    output wire        mb1_FA1_BB0_IO_082_mb1_FB1_BB2_IO_068,
    output wire        mb1_FA1_BB0_IO_083_mb1_FB1_BB2_IO_069,
    output wire        mb1_FA1_BB0_IO_084_mb1_FB1_BB2_IO_086,
    output wire        mb1_FA1_BB0_IO_085_mb1_FB1_BB2_IO_087,
    output wire        mb1_FA1_BB0_IO_086_mb1_FB1_BB2_IO_084,
    output wire        mb1_FA1_BB0_IO_087_mb1_FB1_BB2_IO_085,
    output wire        mb1_FA1_BB0_IO_088_mb1_FB1_BB2_IO_102,
    output wire        mb1_FA1_BB0_IO_089_mb1_FB1_BB2_IO_103,
    output wire        mb1_FA1_BB0_IO_090_mb1_FB1_BB2_IO_080,
    output wire        mb1_FA1_BB0_IO_091_mb1_FB1_BB2_IO_081,
    output wire        mb1_FA1_BB0_IO_092_mb1_FB1_BB2_IO_078,
    output wire        mb1_FA1_BB0_IO_093_mb1_FB1_BB2_IO_079,
    output wire        mb1_FA1_BB0_IO_094_mb1_FB1_BB2_IO_096,
    output wire        mb1_FA1_BB0_IO_095_mb1_FB1_BB2_IO_097,
    output wire        mb1_FA1_BB0_IO_096_mb1_FB1_BB2_IO_094,
    output wire        mb1_FA1_BB0_IO_097_mb1_FB1_BB2_IO_095,
    output wire        mb1_FA1_BB0_IO_098_mb1_FB1_BB2_IO_112,
    output wire        mb1_FA1_BB0_IO_099_mb1_FB1_BB2_IO_113,
    output wire        mb1_FA1_BB0_IO_100_mb1_FB1_BB2_IO_110,
    output wire        mb1_FA1_BB0_IO_101_mb1_FB1_BB2_IO_111,
    output wire        mb1_FA1_BB0_IO_102_mb1_FB1_BB2_IO_088,
    output wire        mb1_FA1_BB0_IO_103_mb1_FB1_BB2_IO_089,
    output wire        mb1_FA1_BB0_IO_104_mb1_FB1_BB2_IO_106,
    output wire        mb1_FA1_BB0_IO_105_mb1_FB1_BB2_IO_107,
    output wire        mb1_FA1_BB0_IO_106_mb1_FB1_BB2_IO_104,
    output wire        mb1_FA1_BB0_IO_107_mb1_FB1_BB2_IO_105,
    output wire        mb1_FA1_BB0_IO_108_mb1_FB1_BB2_IO_122,
    output wire        mb1_FA1_BB0_IO_109_mb1_FB1_BB2_IO_123,
    output wire        mb1_FA1_BB0_IO_110_mb1_FB1_BB2_IO_100,
    output wire        mb1_FA1_BB0_IO_111_mb1_FB1_BB2_IO_101,
    output wire        mb1_FA1_BB0_IO_112_mb1_FB1_BB2_IO_098,
    output wire        mb1_FA1_BB0_IO_113_mb1_FB1_BB2_IO_099,
    output wire        mb1_FA1_BB0_IO_114_mb1_FB1_BB2_IO_116,
    output wire        mb1_FA1_BB0_IO_115_mb1_FB1_BB2_IO_117,
    output wire        mb1_FA1_BB0_IO_116_mb1_FB1_BB2_IO_114,
    output wire        mb1_FA1_BB0_IO_117_mb1_FB1_BB2_IO_115,
    output wire        mb1_FA1_BB0_IO_118_mb1_FB1_BB2_IO_132,
    output wire        mb1_FA1_BB0_IO_119_mb1_FB1_BB2_IO_133,
    output wire        mb1_FA1_BB0_IO_120_mb1_FB1_BB2_IO_130,
    output wire        mb1_FA1_BB0_IO_121_mb1_FB1_BB2_IO_131,
    output wire        mb1_FA1_BB0_IO_122_mb1_FB1_BB2_IO_108,
    output wire        mb1_FA1_BB0_IO_123_mb1_FB1_BB2_IO_109,
    output wire        mb1_FA1_BB0_IO_124_mb1_FB1_BB2_IO_126,
    output wire        mb1_FA1_BB0_IO_125_mb1_FB1_BB2_IO_127,
    output wire        mb1_FA1_BB0_IO_126_mb1_FB1_BB2_IO_124,
    output wire        mb1_FA1_BB0_IO_127_mb1_FB1_BB2_IO_125,
    output wire        mb1_FA1_BB0_IO_130_mb1_FB1_BB2_IO_120,
    output wire        mb1_FA1_BB0_IO_131_mb1_FB1_BB2_IO_121,
    output wire        mb1_FA1_BB0_IO_132_mb1_FB1_BB2_IO_118,
    output wire        mb1_FA1_BB0_IO_133_mb1_FB1_BB2_IO_119,
    output wire        mb1_FA1_BB0_IO_134_mb1_FB1_BB2_IO_136,
    output wire        mb1_FA1_BB0_IO_136_mb1_FB1_BB2_IO_134,
    output wire        mb1_FA1_BB1_CLKIO_N_0_mb1_FA2_BB1_CLKIO_N_7,
    output wire        mb1_FA1_BB1_CLKIO_N_1_mb1_FA2_BB1_CLKIO_N_6,
    output wire        mb1_FA1_BB1_CLKIO_N_2_mb1_FA2_BB1_CLKIO_N_4,
    output wire        mb1_FA1_BB1_CLKIO_N_3_mb1_FA2_BB1_CLKIO_N_3,
    output wire        mb1_FA1_BB1_CLKIO_N_4_mb1_FA2_BB1_CLKIO_N_2,
    output wire        mb1_FA1_BB1_CLKIO_N_5_mb1_FA2_BB1_IO_010,
    output wire        mb1_FA1_BB1_CLKIO_N_6_mb1_FA2_BB1_CLKIO_N_1,
    output wire        mb1_FA1_BB1_CLKIO_N_7_mb1_FA2_BB1_CLKIO_N_0,
    output wire        mb1_FA1_BB1_CLKIO_P_0_mb1_FA2_BB1_CLKIO_P_7,
    output wire        mb1_FA1_BB1_CLKIO_P_1_mb1_FA2_BB1_CLKIO_P_6,
    output wire        mb1_FA1_BB1_CLKIO_P_2_mb1_FA2_BB1_CLKIO_P_4,
    output wire        mb1_FA1_BB1_CLKIO_P_3_mb1_FA2_BB1_CLKIO_P_3,
    output wire        mb1_FA1_BB1_CLKIO_P_4_mb1_FA2_BB1_CLKIO_P_2,
    output wire        mb1_FA1_BB1_CLKIO_P_5_mb1_FA2_BB1_IO_011,
    output wire        mb1_FA1_BB1_CLKIO_P_6_mb1_FA2_BB1_CLKIO_P_1,
    output wire        mb1_FA1_BB1_CLKIO_P_7_mb1_FA2_BB1_CLKIO_P_0,
    output wire        mb1_FA1_BB1_IO_004_mb1_FA2_BB1_IO_006,
    output wire        mb1_FA1_BB1_IO_005_mb1_FA2_BB1_IO_007,
    output wire        mb1_FA1_BB1_IO_006_mb1_FA2_BB1_IO_004,
    output wire        mb1_FA1_BB1_IO_007_mb1_FA2_BB1_IO_005,
    output wire        mb1_FA1_BB1_IO_008_mb1_FA2_BB1_IO_022,
    output wire        mb1_FA1_BB1_IO_009_mb1_FA2_BB1_IO_023,
    output wire        mb1_FA1_BB1_IO_010_mb1_FA2_BB1_CLKIO_N_5,
    output wire        mb1_FA1_BB1_IO_011_mb1_FA2_BB1_CLKIO_P_5,
    output wire        mb1_FA1_BB1_IO_012_mb1_FA2_BB1_IO_012,
    output wire        mb1_FA1_BB1_IO_013_mb1_FA2_BB1_IO_013,
    output wire        mb1_FA1_BB1_IO_014_mb1_FA2_BB1_IO_016,
    output wire        mb1_FA1_BB1_IO_015_mb1_FA2_BB1_IO_017,
    output wire        mb1_FA1_BB1_IO_016_mb1_FA2_BB1_IO_014,
    output wire        mb1_FA1_BB1_IO_017_mb1_FA2_BB1_IO_015,
    output wire        mb1_FA1_BB1_IO_018_mb1_FA2_BB1_IO_032,
    output wire        mb1_FA1_BB1_IO_019_mb1_FA2_BB1_IO_033,
    output wire        mb1_FA1_BB1_IO_020_mb1_FA2_BB1_IO_030,
    output wire        mb1_FA1_BB1_IO_021_mb1_FA2_BB1_IO_031,
    output wire        mb1_FA1_BB1_IO_022_mb1_FA2_BB1_IO_008,
    output wire        mb1_FA1_BB1_IO_023_mb1_FA2_BB1_IO_009,
    output wire        mb1_FA1_BB1_IO_024_mb1_FA2_BB1_IO_026,
    output wire        mb1_FA1_BB1_IO_025_mb1_FA2_BB1_IO_027,
    output wire        mb1_FA1_BB1_IO_026_mb1_FA2_BB1_IO_024,
    output wire        mb1_FA1_BB1_IO_027_mb1_FA2_BB1_IO_025,
    output wire        mb1_FA1_BB1_IO_028_mb1_FA2_BB1_IO_042,
    output wire        mb1_FA1_BB1_IO_029_mb1_FA2_BB1_IO_043,
    output wire        mb1_FA1_BB1_IO_030_mb1_FA2_BB1_IO_020,
    output wire        mb1_FA1_BB1_IO_031_mb1_FA2_BB1_IO_021,
    output wire        mb1_FA1_BB1_IO_032_mb1_FA2_BB1_IO_018,
    output wire        mb1_FA1_BB1_IO_033_mb1_FA2_BB1_IO_019,
    output wire        mb1_FA1_BB1_IO_034_mb1_FA2_BB1_IO_036,
    output wire        mb1_FA1_BB1_IO_035_mb1_FA2_BB1_IO_037,
    output wire        mb1_FA1_BB1_IO_036_mb1_FA2_BB1_IO_034,
    output wire        mb1_FA1_BB1_IO_037_mb1_FA2_BB1_IO_035,
    output wire        mb1_FA1_BB1_IO_038_mb1_FA2_BB1_IO_052,
    output wire        mb1_FA1_BB1_IO_039_mb1_FA2_BB1_IO_053,
    output wire        mb1_FA1_BB1_IO_040_mb1_FA2_BB1_IO_050,
    output wire        mb1_FA1_BB1_IO_041_mb1_FA2_BB1_IO_051,
    output wire        mb1_FA1_BB1_IO_042_mb1_FA2_BB1_IO_028,
    output wire        mb1_FA1_BB1_IO_043_mb1_FA2_BB1_IO_029,
    output wire        mb1_FA1_BB1_IO_044_mb1_FA2_BB1_IO_046,
    output wire        mb1_FA1_BB1_IO_045_mb1_FA2_BB1_IO_047,
    output wire        mb1_FA1_BB1_IO_046_mb1_FA2_BB1_IO_044,
    output wire        mb1_FA1_BB1_IO_047_mb1_FA2_BB1_IO_045,
    output wire        mb1_FA1_BB1_IO_048_mb1_FA2_BB1_IO_062,
    output wire        mb1_FA1_BB1_IO_049_mb1_FA2_BB1_IO_063,
    output wire        mb1_FA1_BB1_IO_050_mb1_FA2_BB1_IO_040,
    output wire        mb1_FA1_BB1_IO_051_mb1_FA2_BB1_IO_041,
    output wire        mb1_FA1_BB1_IO_052_mb1_FA2_BB1_IO_038,
    output wire        mb1_FA1_BB1_IO_053_mb1_FA2_BB1_IO_039,
    output wire        mb1_FA1_BB1_IO_054_mb1_FA2_BB1_IO_056,
    output wire        mb1_FA1_BB1_IO_055_mb1_FA2_BB1_IO_057,
    output wire        mb1_FA1_BB1_IO_056_mb1_FA2_BB1_IO_054,
    output wire        mb1_FA1_BB1_IO_057_mb1_FA2_BB1_IO_055,
    output wire        mb1_FA1_BB1_IO_058_mb1_FA2_BB1_IO_072,
    output wire        mb1_FA1_BB1_IO_059_mb1_FA2_BB1_IO_073,
    output wire        mb1_FA1_BB1_IO_060_mb1_FA2_BB1_IO_070,
    output wire        mb1_FA1_BB1_IO_061_mb1_FA2_BB1_IO_071,
    output wire        mb1_FA1_BB1_IO_062_mb1_FA2_BB1_IO_048,
    output wire        mb1_FA1_BB1_IO_063_mb1_FA2_BB1_IO_049,
    output wire        mb1_FA1_BB1_IO_064_mb1_FA2_BB1_IO_066,
    output wire        mb1_FA1_BB1_IO_065_mb1_FA2_BB1_IO_067,
    output wire        mb1_FA1_BB1_IO_066_mb1_FA2_BB1_IO_064,
    output wire        mb1_FA1_BB1_IO_067_mb1_FA2_BB1_IO_065,
    output wire        mb1_FA1_BB1_IO_068_mb1_FA2_BB1_IO_082,
    output wire        mb1_FA1_BB1_IO_069_mb1_FA2_BB1_IO_083,
    output wire        mb1_FA1_BB1_IO_070_mb1_FA2_BB1_IO_060,
    output wire        mb1_FA1_BB1_IO_071_mb1_FA2_BB1_IO_061,
    output wire        mb1_FA1_BB1_IO_072_mb1_FA2_BB1_IO_058,
    output wire        mb1_FA1_BB1_IO_073_mb1_FA2_BB1_IO_059,
    output wire        mb1_FA1_BB1_IO_074_mb1_FA2_BB1_IO_076,
    output wire        mb1_FA1_BB1_IO_075_mb1_FA2_BB1_IO_077,
    output wire        mb1_FA1_BB1_IO_076_mb1_FA2_BB1_IO_074,
    output wire        mb1_FA1_BB1_IO_077_mb1_FA2_BB1_IO_075,
    output wire        mb1_FA1_BB1_IO_078_mb1_FA2_BB1_IO_092,
    output wire        mb1_FA1_BB1_IO_079_mb1_FA2_BB1_IO_093,
    output wire        mb1_FA1_BB1_IO_080_mb1_FA2_BB1_IO_090,
    output wire        mb1_FA1_BB1_IO_081_mb1_FA2_BB1_IO_091,
    output wire        mb1_FA1_BB1_IO_082_mb1_FA2_BB1_IO_068,
    output wire        mb1_FA1_BB1_IO_083_mb1_FA2_BB1_IO_069,
    output wire        mb1_FA1_BB1_IO_084_mb1_FA2_BB1_IO_086,
    output wire        mb1_FA1_BB1_IO_085_mb1_FA2_BB1_IO_087,
    output wire        mb1_FA1_BB1_IO_086_mb1_FA2_BB1_IO_084,
    output wire        mb1_FA1_BB1_IO_087_mb1_FA2_BB1_IO_085,
    output wire        mb1_FA1_BB1_IO_088_mb1_FA2_BB1_IO_102,
    output wire        mb1_FA1_BB1_IO_089_mb1_FA2_BB1_IO_103,
    output wire        mb1_FA1_BB1_IO_090_mb1_FA2_BB1_IO_080,
    output wire        mb1_FA1_BB1_IO_091_mb1_FA2_BB1_IO_081,
    output wire        mb1_FA1_BB1_IO_092_mb1_FA2_BB1_IO_078,
    output wire        mb1_FA1_BB1_IO_093_mb1_FA2_BB1_IO_079,
    output wire        mb1_FA1_BB1_IO_094_mb1_FA2_BB1_IO_096,
    output wire        mb1_FA1_BB1_IO_095_mb1_FA2_BB1_IO_097,
    output wire        mb1_FA1_BB1_IO_096_mb1_FA2_BB1_IO_094,
    output wire        mb1_FA1_BB1_IO_097_mb1_FA2_BB1_IO_095,
    output wire        mb1_FA1_BB1_IO_098_mb1_FA2_BB1_IO_112,
    output wire        mb1_FA1_BB1_IO_099_mb1_FA2_BB1_IO_113,
    output wire        mb1_FA1_BB1_IO_100_mb1_FA2_BB1_IO_110,
    output wire        mb1_FA1_BB1_IO_101_mb1_FA2_BB1_IO_111,
    output wire        mb1_FA1_BB1_IO_102_mb1_FA2_BB1_IO_088,
    output wire        mb1_FA1_BB1_IO_103_mb1_FA2_BB1_IO_089,
    output wire        mb1_FA1_BB1_IO_104_mb1_FA2_BB1_IO_106,
    output wire        mb1_FA1_BB1_IO_105_mb1_FA2_BB1_IO_107,
    output wire        mb1_FA1_BB1_IO_106_mb1_FA2_BB1_IO_104,
    output wire        mb1_FA1_BB1_IO_107_mb1_FA2_BB1_IO_105,
    output wire        mb1_FA1_BB1_IO_108_mb1_FA2_BB1_IO_122,
    output wire        mb1_FA1_BB1_IO_109_mb1_FA2_BB1_IO_123,
    output wire        mb1_FA1_BB1_IO_110_mb1_FA2_BB1_IO_100,
    output wire        mb1_FA1_BB1_IO_111_mb1_FA2_BB1_IO_101,
    output wire        mb1_FA1_BB1_IO_112_mb1_FA2_BB1_IO_098,
    output wire        mb1_FA1_BB1_IO_113_mb1_FA2_BB1_IO_099,
    output wire        mb1_FA1_BB1_IO_114_mb1_FA2_BB1_IO_116,
    output wire        mb1_FA1_BB1_IO_115_mb1_FA2_BB1_IO_117,
    output wire        mb1_FA1_BB1_IO_116_mb1_FA2_BB1_IO_114,
    output wire        mb1_FA1_BB1_IO_117_mb1_FA2_BB1_IO_115,
    output wire        mb1_FA1_BB1_IO_118_mb1_FA2_BB1_IO_132,
    output wire        mb1_FA1_BB1_IO_119_mb1_FA2_BB1_IO_133,
    output wire        mb1_FA1_BB1_IO_120_mb1_FA2_BB1_IO_130,
    output wire        mb1_FA1_BB1_IO_121_mb1_FA2_BB1_IO_131,
    output wire        mb1_FA1_BB1_IO_122_mb1_FA2_BB1_IO_108,
    output wire        mb1_FA1_BB1_IO_123_mb1_FA2_BB1_IO_109,
    output wire        mb1_FA1_BB1_IO_124_mb1_FA2_BB1_IO_126,
    output wire        mb1_FA1_BB1_IO_125_mb1_FA2_BB1_IO_127,
    output wire        mb1_FA1_BB1_IO_126_mb1_FA2_BB1_IO_124,
    output wire        mb1_FA1_BB1_IO_127_mb1_FA2_BB1_IO_125,
    output wire        mb1_FA1_BB1_IO_130_mb1_FA2_BB1_IO_120,
    output wire        mb1_FA1_BB1_IO_131_mb1_FA2_BB1_IO_121,
    output wire        mb1_FA1_BB1_IO_132_mb1_FA2_BB1_IO_118,
    output wire        mb1_FA1_BB1_IO_133_mb1_FA2_BB1_IO_119,
    output wire        mb1_FA1_BB1_IO_134_mb1_FA2_BB1_IO_136,
    output wire        mb1_FA1_BB1_IO_136_mb1_FA2_BB1_IO_134);

  localparam TX_PINS            = 1314;
  localparam RX_PINS            = 0;
  localparam USE_CLK_INPUT_BUFG = 0;

  wire [TX_PINS-1:0] tx_pin;

  assign mb1_FA1_TA1_CLKIO_N_0_mb1_FB1_TA2_CLKIO_N_7 = tx_pin[0];
  assign mb1_FA1_TA1_CLKIO_N_1_mb1_FB1_TA2_CLKIO_N_6 = tx_pin[1];
  assign mb1_FA1_TA1_CLKIO_N_2_mb1_FB1_TA2_CLKIO_N_4 = tx_pin[2];
  assign mb1_FA1_TA1_CLKIO_N_3_mb1_FB1_TA2_CLKIO_N_3 = tx_pin[3];
  assign mb1_FA1_TA1_CLKIO_N_4_mb1_FB1_TA2_CLKIO_N_2 = tx_pin[4];
  assign mb1_FA1_TA1_CLKIO_N_5_mb1_FB1_TA2_IO_010 = tx_pin[5];
  assign mb1_FA1_TA1_CLKIO_N_6_mb1_FB1_TA2_CLKIO_N_1 = tx_pin[6];
  assign mb1_FA1_TA1_CLKIO_N_7_mb1_FB1_TA2_CLKIO_N_0 = tx_pin[7];
  assign mb1_FA1_TA1_CLKIO_P_0_mb1_FB1_TA2_CLKIO_P_7 = tx_pin[8];
  assign mb1_FA1_TA1_CLKIO_P_1_mb1_FB1_TA2_CLKIO_P_6 = tx_pin[9];
  assign mb1_FA1_TA1_CLKIO_P_2_mb1_FB1_TA2_CLKIO_P_4 = tx_pin[10];
  assign mb1_FA1_TA1_CLKIO_P_3_mb1_FB1_TA2_CLKIO_P_3 = tx_pin[11];
  assign mb1_FA1_TA1_CLKIO_P_4_mb1_FB1_TA2_CLKIO_P_2 = tx_pin[12];
  assign mb1_FA1_TA1_CLKIO_P_5_mb1_FB1_TA2_IO_011 = tx_pin[13];
  assign mb1_FA1_TA1_CLKIO_P_6_mb1_FB1_TA2_CLKIO_P_1 = tx_pin[14];
  assign mb1_FA1_TA1_CLKIO_P_7_mb1_FB1_TA2_CLKIO_P_0 = tx_pin[15];
  assign mb1_FA1_TA1_IO_004_mb1_FB1_TA2_IO_006 = tx_pin[16];
  assign mb1_FA1_TA1_IO_005_mb1_FB1_TA2_IO_007 = tx_pin[17];
  assign mb1_FA1_TA1_IO_006_mb1_FB1_TA2_IO_004 = tx_pin[18];
  assign mb1_FA1_TA1_IO_007_mb1_FB1_TA2_IO_005 = tx_pin[19];
  assign mb1_FA1_TA1_IO_008_mb1_FB1_TA2_IO_022 = tx_pin[20];
  assign mb1_FA1_TA1_IO_009_mb1_FB1_TA2_IO_023 = tx_pin[21];
  assign mb1_FA1_TA1_IO_010_mb1_FB1_TA2_CLKIO_N_5 = tx_pin[22];
  assign mb1_FA1_TA1_IO_011_mb1_FB1_TA2_CLKIO_P_5 = tx_pin[23];
  assign mb1_FA1_TA1_IO_012_mb1_FB1_TA2_IO_012 = tx_pin[24];
  assign mb1_FA1_TA1_IO_013_mb1_FB1_TA2_IO_013 = tx_pin[25];
  assign mb1_FA1_TA1_IO_014_mb1_FB1_TA2_IO_016 = tx_pin[26];
  assign mb1_FA1_TA1_IO_015_mb1_FB1_TA2_IO_017 = tx_pin[27];
  assign mb1_FA1_TA1_IO_016_mb1_FB1_TA2_IO_014 = tx_pin[28];
  assign mb1_FA1_TA1_IO_017_mb1_FB1_TA2_IO_015 = tx_pin[29];
  assign mb1_FA1_TA1_IO_018_mb1_FB1_TA2_IO_032 = tx_pin[30];
  assign mb1_FA1_TA1_IO_019_mb1_FB1_TA2_IO_033 = tx_pin[31];
  assign mb1_FA1_TA1_IO_020_mb1_FB1_TA2_IO_030 = tx_pin[32];
  assign mb1_FA1_TA1_IO_021_mb1_FB1_TA2_IO_031 = tx_pin[33];
  assign mb1_FA1_TA1_IO_022_mb1_FB1_TA2_IO_008 = tx_pin[34];
  assign mb1_FA1_TA1_IO_023_mb1_FB1_TA2_IO_009 = tx_pin[35];
  assign mb1_FA1_TA1_IO_024_mb1_FB1_TA2_IO_026 = tx_pin[36];
  assign mb1_FA1_TA1_IO_025_mb1_FB1_TA2_IO_027 = tx_pin[37];
  assign mb1_FA1_TA1_IO_026_mb1_FB1_TA2_IO_024 = tx_pin[38];
  assign mb1_FA1_TA1_IO_027_mb1_FB1_TA2_IO_025 = tx_pin[39];
  assign mb1_FA1_TA1_IO_028_mb1_FB1_TA2_IO_042 = tx_pin[40];
  assign mb1_FA1_TA1_IO_029_mb1_FB1_TA2_IO_043 = tx_pin[41];
  assign mb1_FA1_TA1_IO_030_mb1_FB1_TA2_IO_020 = tx_pin[42];
  assign mb1_FA1_TA1_IO_031_mb1_FB1_TA2_IO_021 = tx_pin[43];
  assign mb1_FA1_TA1_IO_032_mb1_FB1_TA2_IO_018 = tx_pin[44];
  assign mb1_FA1_TA1_IO_033_mb1_FB1_TA2_IO_019 = tx_pin[45];
  assign mb1_FA1_TA1_IO_034_mb1_FB1_TA2_IO_036 = tx_pin[46];
  assign mb1_FA1_TA1_IO_035_mb1_FB1_TA2_IO_037 = tx_pin[47];
  assign mb1_FA1_TA1_IO_036_mb1_FB1_TA2_IO_034 = tx_pin[48];
  assign mb1_FA1_TA1_IO_037_mb1_FB1_TA2_IO_035 = tx_pin[49];
  assign mb1_FA1_TA1_IO_038_mb1_FB1_TA2_IO_052 = tx_pin[50];
  assign mb1_FA1_TA1_IO_039_mb1_FB1_TA2_IO_053 = tx_pin[51];
  assign mb1_FA1_TA1_IO_040_mb1_FB1_TA2_IO_050 = tx_pin[52];
  assign mb1_FA1_TA1_IO_041_mb1_FB1_TA2_IO_051 = tx_pin[53];
  assign mb1_FA1_TA1_IO_042_mb1_FB1_TA2_IO_028 = tx_pin[54];
  assign mb1_FA1_TA1_IO_043_mb1_FB1_TA2_IO_029 = tx_pin[55];
  assign mb1_FA1_TA1_IO_044_mb1_FB1_TA2_IO_046 = tx_pin[56];
  assign mb1_FA1_TA1_IO_045_mb1_FB1_TA2_IO_047 = tx_pin[57];
  assign mb1_FA1_TA1_IO_046_mb1_FB1_TA2_IO_044 = tx_pin[58];
  assign mb1_FA1_TA1_IO_047_mb1_FB1_TA2_IO_045 = tx_pin[59];
  assign mb1_FA1_TA1_IO_048_mb1_FB1_TA2_IO_062 = tx_pin[60];
  assign mb1_FA1_TA1_IO_049_mb1_FB1_TA2_IO_063 = tx_pin[61];
  assign mb1_FA1_TA1_IO_050_mb1_FB1_TA2_IO_040 = tx_pin[62];
  assign mb1_FA1_TA1_IO_051_mb1_FB1_TA2_IO_041 = tx_pin[63];
  assign mb1_FA1_TA1_IO_052_mb1_FB1_TA2_IO_038 = tx_pin[64];
  assign mb1_FA1_TA1_IO_053_mb1_FB1_TA2_IO_039 = tx_pin[65];
  assign mb1_FA1_TA1_IO_054_mb1_FB1_TA2_IO_056 = tx_pin[66];
  assign mb1_FA1_TA1_IO_055_mb1_FB1_TA2_IO_057 = tx_pin[67];
  assign mb1_FA1_TA1_IO_056_mb1_FB1_TA2_IO_054 = tx_pin[68];
  assign mb1_FA1_TA1_IO_057_mb1_FB1_TA2_IO_055 = tx_pin[69];
  assign mb1_FA1_TA1_IO_058_mb1_FB1_TA2_IO_072 = tx_pin[70];
  assign mb1_FA1_TA1_IO_059_mb1_FB1_TA2_IO_073 = tx_pin[71];
  assign mb1_FA1_TA1_IO_060_mb1_FB1_TA2_IO_070 = tx_pin[72];
  assign mb1_FA1_TA1_IO_061_mb1_FB1_TA2_IO_071 = tx_pin[73];
  assign mb1_FA1_TA1_IO_062_mb1_FB1_TA2_IO_048 = tx_pin[74];
  assign mb1_FA1_TA1_IO_063_mb1_FB1_TA2_IO_049 = tx_pin[75];
  assign mb1_FA1_TA1_IO_064_mb1_FB1_TA2_IO_066 = tx_pin[76];
  assign mb1_FA1_TA1_IO_065_mb1_FB1_TA2_IO_067 = tx_pin[77];
  assign mb1_FA1_TA1_IO_066_mb1_FB1_TA2_IO_064 = tx_pin[78];
  assign mb1_FA1_TA1_IO_067_mb1_FB1_TA2_IO_065 = tx_pin[79];
  assign mb1_FA1_TA1_IO_068_mb1_FB1_TA2_IO_082 = tx_pin[80];
  assign mb1_FA1_TA1_IO_069_mb1_FB1_TA2_IO_083 = tx_pin[81];
  assign mb1_FA1_TA1_IO_070_mb1_FB1_TA2_IO_060 = tx_pin[82];
  assign mb1_FA1_TA1_IO_071_mb1_FB1_TA2_IO_061 = tx_pin[83];
  assign mb1_FA1_TA1_IO_072_mb1_FB1_TA2_IO_058 = tx_pin[84];
  assign mb1_FA1_TA1_IO_073_mb1_FB1_TA2_IO_059 = tx_pin[85];
  assign mb1_FA1_TA1_IO_074_mb1_FB1_TA2_IO_076 = tx_pin[86];
  assign mb1_FA1_TA1_IO_075_mb1_FB1_TA2_IO_077 = tx_pin[87];
  assign mb1_FA1_TA1_IO_076_mb1_FB1_TA2_IO_074 = tx_pin[88];
  assign mb1_FA1_TA1_IO_077_mb1_FB1_TA2_IO_075 = tx_pin[89];
  assign mb1_FA1_TA1_IO_078_mb1_FB1_TA2_IO_092 = tx_pin[90];
  assign mb1_FA1_TA1_IO_079_mb1_FB1_TA2_IO_093 = tx_pin[91];
  assign mb1_FA1_TA1_IO_080_mb1_FB1_TA2_IO_090 = tx_pin[92];
  assign mb1_FA1_TA1_IO_081_mb1_FB1_TA2_IO_091 = tx_pin[93];
  assign mb1_FA1_TA1_IO_082_mb1_FB1_TA2_IO_068 = tx_pin[94];
  assign mb1_FA1_TA1_IO_083_mb1_FB1_TA2_IO_069 = tx_pin[95];
  assign mb1_FA1_TA1_IO_084_mb1_FB1_TA2_IO_086 = tx_pin[96];
  assign mb1_FA1_TA1_IO_085_mb1_FB1_TA2_IO_087 = tx_pin[97];
  assign mb1_FA1_TA1_IO_086_mb1_FB1_TA2_IO_084 = tx_pin[98];
  assign mb1_FA1_TA1_IO_087_mb1_FB1_TA2_IO_085 = tx_pin[99];
  assign mb1_FA1_TA1_IO_088_mb1_FB1_TA2_IO_102 = tx_pin[100];
  assign mb1_FA1_TA1_IO_089_mb1_FB1_TA2_IO_103 = tx_pin[101];
  assign mb1_FA1_TA1_IO_090_mb1_FB1_TA2_IO_080 = tx_pin[102];
  assign mb1_FA1_TA1_IO_091_mb1_FB1_TA2_IO_081 = tx_pin[103];
  assign mb1_FA1_TA1_IO_092_mb1_FB1_TA2_IO_078 = tx_pin[104];
  assign mb1_FA1_TA1_IO_093_mb1_FB1_TA2_IO_079 = tx_pin[105];
  assign mb1_FA1_TA1_IO_094_mb1_FB1_TA2_IO_096 = tx_pin[106];
  assign mb1_FA1_TA1_IO_095_mb1_FB1_TA2_IO_097 = tx_pin[107];
  assign mb1_FA1_TA1_IO_096_mb1_FB1_TA2_IO_094 = tx_pin[108];
  assign mb1_FA1_TA1_IO_097_mb1_FB1_TA2_IO_095 = tx_pin[109];
  assign mb1_FA1_TA1_IO_098_mb1_FB1_TA2_IO_112 = tx_pin[110];
  assign mb1_FA1_TA1_IO_099_mb1_FB1_TA2_IO_113 = tx_pin[111];
  assign mb1_FA1_TA1_IO_100_mb1_FB1_TA2_IO_110 = tx_pin[112];
  assign mb1_FA1_TA1_IO_101_mb1_FB1_TA2_IO_111 = tx_pin[113];
  assign mb1_FA1_TA1_IO_102_mb1_FB1_TA2_IO_088 = tx_pin[114];
  assign mb1_FA1_TA1_IO_103_mb1_FB1_TA2_IO_089 = tx_pin[115];
  assign mb1_FA1_TA1_IO_104_mb1_FB1_TA2_IO_106 = tx_pin[116];
  assign mb1_FA1_TA1_IO_105_mb1_FB1_TA2_IO_107 = tx_pin[117];
  assign mb1_FA1_TA1_IO_106_mb1_FB1_TA2_IO_104 = tx_pin[118];
  assign mb1_FA1_TA1_IO_107_mb1_FB1_TA2_IO_105 = tx_pin[119];
  assign mb1_FA1_TA1_IO_108_mb1_FB1_TA2_IO_122 = tx_pin[120];
  assign mb1_FA1_TA1_IO_109_mb1_FB1_TA2_IO_123 = tx_pin[121];
  assign mb1_FA1_TA1_IO_110_mb1_FB1_TA2_IO_100 = tx_pin[122];
  assign mb1_FA1_TA1_IO_111_mb1_FB1_TA2_IO_101 = tx_pin[123];
  assign mb1_FA1_TA1_IO_112_mb1_FB1_TA2_IO_098 = tx_pin[124];
  assign mb1_FA1_TA1_IO_113_mb1_FB1_TA2_IO_099 = tx_pin[125];
  assign mb1_FA1_TA1_IO_114_mb1_FB1_TA2_IO_116 = tx_pin[126];
  assign mb1_FA1_TA1_IO_115_mb1_FB1_TA2_IO_117 = tx_pin[127];
  assign mb1_FA1_TA1_IO_116_mb1_FB1_TA2_IO_114 = tx_pin[128];
  assign mb1_FA1_TA1_IO_117_mb1_FB1_TA2_IO_115 = tx_pin[129];
  assign mb1_FA1_TA1_IO_118_mb1_FB1_TA2_IO_132 = tx_pin[130];
  assign mb1_FA1_TA1_IO_119_mb1_FB1_TA2_IO_133 = tx_pin[131];
  assign mb1_FA1_TA1_IO_120_mb1_FB1_TA2_IO_130 = tx_pin[132];
  assign mb1_FA1_TA1_IO_121_mb1_FB1_TA2_IO_131 = tx_pin[133];
  assign mb1_FA1_TA1_IO_122_mb1_FB1_TA2_IO_108 = tx_pin[134];
  assign mb1_FA1_TA1_IO_123_mb1_FB1_TA2_IO_109 = tx_pin[135];
  assign mb1_FA1_TA1_IO_124_mb1_FB1_TA2_IO_126 = tx_pin[136];
  assign mb1_FA1_TA1_IO_125_mb1_FB1_TA2_IO_127 = tx_pin[137];
  assign mb1_FA1_TA1_IO_126_mb1_FB1_TA2_IO_124 = tx_pin[138];
  assign mb1_FA1_TA1_IO_127_mb1_FB1_TA2_IO_125 = tx_pin[139];
  assign mb1_FA1_TA1_IO_130_mb1_FB1_TA2_IO_120 = tx_pin[140];
  assign mb1_FA1_TA1_IO_131_mb1_FB1_TA2_IO_121 = tx_pin[141];
  assign mb1_FA1_TA1_IO_132_mb1_FB1_TA2_IO_118 = tx_pin[142];
  assign mb1_FA1_TA1_IO_133_mb1_FB1_TA2_IO_119 = tx_pin[143];
  assign mb1_FA1_TA1_IO_134_mb1_FB1_TA2_IO_136 = tx_pin[144];
  assign mb1_FA1_TA1_IO_136_mb1_FB1_TA2_IO_134 = tx_pin[145];
  assign mb1_FA1_TB0_CLKIO_N_0_mb1_FB1_TB2_CLKIO_N_7 = tx_pin[146];
  assign mb1_FA1_TB0_CLKIO_N_1_mb1_FB1_TB2_CLKIO_N_6 = tx_pin[147];
  assign mb1_FA1_TB0_CLKIO_N_2_mb1_FB1_TB2_CLKIO_N_4 = tx_pin[148];
  assign mb1_FA1_TB0_CLKIO_N_3_mb1_FB1_TB2_CLKIO_N_3 = tx_pin[149];
  assign mb1_FA1_TB0_CLKIO_N_4_mb1_FB1_TB2_CLKIO_N_2 = tx_pin[150];
  assign mb1_FA1_TB0_CLKIO_N_5_mb1_FB1_TB2_IO_010 = tx_pin[151];
  assign mb1_FA1_TB0_CLKIO_N_6_mb1_FB1_TB2_CLKIO_N_1 = tx_pin[152];
  assign mb1_FA1_TB0_CLKIO_N_7_mb1_FB1_TB2_CLKIO_N_0 = tx_pin[153];
  assign mb1_FA1_TB0_CLKIO_P_0_mb1_FB1_TB2_CLKIO_P_7 = tx_pin[154];
  assign mb1_FA1_TB0_CLKIO_P_1_mb1_FB1_TB2_CLKIO_P_6 = tx_pin[155];
  assign mb1_FA1_TB0_CLKIO_P_2_mb1_FB1_TB2_CLKIO_P_4 = tx_pin[156];
  assign mb1_FA1_TB0_CLKIO_P_3_mb1_FB1_TB2_CLKIO_P_3 = tx_pin[157];
  assign mb1_FA1_TB0_CLKIO_P_4_mb1_FB1_TB2_CLKIO_P_2 = tx_pin[158];
  assign mb1_FA1_TB0_CLKIO_P_5_mb1_FB1_TB2_IO_011 = tx_pin[159];
  assign mb1_FA1_TB0_CLKIO_P_6_mb1_FB1_TB2_CLKIO_P_1 = tx_pin[160];
  assign mb1_FA1_TB0_CLKIO_P_7_mb1_FB1_TB2_CLKIO_P_0 = tx_pin[161];
  assign mb1_FA1_TB0_IO_004_mb1_FB1_TB2_IO_006 = tx_pin[162];
  assign mb1_FA1_TB0_IO_005_mb1_FB1_TB2_IO_007 = tx_pin[163];
  assign mb1_FA1_TB0_IO_006_mb1_FB1_TB2_IO_004 = tx_pin[164];
  assign mb1_FA1_TB0_IO_007_mb1_FB1_TB2_IO_005 = tx_pin[165];
  assign mb1_FA1_TB0_IO_008_mb1_FB1_TB2_IO_022 = tx_pin[166];
  assign mb1_FA1_TB0_IO_009_mb1_FB1_TB2_IO_023 = tx_pin[167];
  assign mb1_FA1_TB0_IO_010_mb1_FB1_TB2_CLKIO_N_5 = tx_pin[168];
  assign mb1_FA1_TB0_IO_011_mb1_FB1_TB2_CLKIO_P_5 = tx_pin[169];
  assign mb1_FA1_TB0_IO_012_mb1_FB1_TB2_IO_012 = tx_pin[170];
  assign mb1_FA1_TB0_IO_013_mb1_FB1_TB2_IO_013 = tx_pin[171];
  assign mb1_FA1_TB0_IO_014_mb1_FB1_TB2_IO_016 = tx_pin[172];
  assign mb1_FA1_TB0_IO_015_mb1_FB1_TB2_IO_017 = tx_pin[173];
  assign mb1_FA1_TB0_IO_016_mb1_FB1_TB2_IO_014 = tx_pin[174];
  assign mb1_FA1_TB0_IO_017_mb1_FB1_TB2_IO_015 = tx_pin[175];
  assign mb1_FA1_TB0_IO_018_mb1_FB1_TB2_IO_032 = tx_pin[176];
  assign mb1_FA1_TB0_IO_019_mb1_FB1_TB2_IO_033 = tx_pin[177];
  assign mb1_FA1_TB0_IO_020_mb1_FB1_TB2_IO_030 = tx_pin[178];
  assign mb1_FA1_TB0_IO_021_mb1_FB1_TB2_IO_031 = tx_pin[179];
  assign mb1_FA1_TB0_IO_022_mb1_FB1_TB2_IO_008 = tx_pin[180];
  assign mb1_FA1_TB0_IO_023_mb1_FB1_TB2_IO_009 = tx_pin[181];
  assign mb1_FA1_TB0_IO_024_mb1_FB1_TB2_IO_026 = tx_pin[182];
  assign mb1_FA1_TB0_IO_025_mb1_FB1_TB2_IO_027 = tx_pin[183];
  assign mb1_FA1_TB0_IO_026_mb1_FB1_TB2_IO_024 = tx_pin[184];
  assign mb1_FA1_TB0_IO_027_mb1_FB1_TB2_IO_025 = tx_pin[185];
  assign mb1_FA1_TB0_IO_028_mb1_FB1_TB2_IO_042 = tx_pin[186];
  assign mb1_FA1_TB0_IO_029_mb1_FB1_TB2_IO_043 = tx_pin[187];
  assign mb1_FA1_TB0_IO_030_mb1_FB1_TB2_IO_020 = tx_pin[188];
  assign mb1_FA1_TB0_IO_031_mb1_FB1_TB2_IO_021 = tx_pin[189];
  assign mb1_FA1_TB0_IO_032_mb1_FB1_TB2_IO_018 = tx_pin[190];
  assign mb1_FA1_TB0_IO_033_mb1_FB1_TB2_IO_019 = tx_pin[191];
  assign mb1_FA1_TB0_IO_034_mb1_FB1_TB2_IO_036 = tx_pin[192];
  assign mb1_FA1_TB0_IO_035_mb1_FB1_TB2_IO_037 = tx_pin[193];
  assign mb1_FA1_TB0_IO_036_mb1_FB1_TB2_IO_034 = tx_pin[194];
  assign mb1_FA1_TB0_IO_037_mb1_FB1_TB2_IO_035 = tx_pin[195];
  assign mb1_FA1_TB0_IO_038_mb1_FB1_TB2_IO_052 = tx_pin[196];
  assign mb1_FA1_TB0_IO_039_mb1_FB1_TB2_IO_053 = tx_pin[197];
  assign mb1_FA1_TB0_IO_040_mb1_FB1_TB2_IO_050 = tx_pin[198];
  assign mb1_FA1_TB0_IO_041_mb1_FB1_TB2_IO_051 = tx_pin[199];
  assign mb1_FA1_TB0_IO_042_mb1_FB1_TB2_IO_028 = tx_pin[200];
  assign mb1_FA1_TB0_IO_043_mb1_FB1_TB2_IO_029 = tx_pin[201];
  assign mb1_FA1_TB0_IO_044_mb1_FB1_TB2_IO_046 = tx_pin[202];
  assign mb1_FA1_TB0_IO_045_mb1_FB1_TB2_IO_047 = tx_pin[203];
  assign mb1_FA1_TB0_IO_046_mb1_FB1_TB2_IO_044 = tx_pin[204];
  assign mb1_FA1_TB0_IO_047_mb1_FB1_TB2_IO_045 = tx_pin[205];
  assign mb1_FA1_TB0_IO_048_mb1_FB1_TB2_IO_062 = tx_pin[206];
  assign mb1_FA1_TB0_IO_049_mb1_FB1_TB2_IO_063 = tx_pin[207];
  assign mb1_FA1_TB0_IO_050_mb1_FB1_TB2_IO_040 = tx_pin[208];
  assign mb1_FA1_TB0_IO_051_mb1_FB1_TB2_IO_041 = tx_pin[209];
  assign mb1_FA1_TB0_IO_052_mb1_FB1_TB2_IO_038 = tx_pin[210];
  assign mb1_FA1_TB0_IO_053_mb1_FB1_TB2_IO_039 = tx_pin[211];
  assign mb1_FA1_TB0_IO_054_mb1_FB1_TB2_IO_056 = tx_pin[212];
  assign mb1_FA1_TB0_IO_055_mb1_FB1_TB2_IO_057 = tx_pin[213];
  assign mb1_FA1_TB0_IO_056_mb1_FB1_TB2_IO_054 = tx_pin[214];
  assign mb1_FA1_TB0_IO_057_mb1_FB1_TB2_IO_055 = tx_pin[215];
  assign mb1_FA1_TB0_IO_058_mb1_FB1_TB2_IO_072 = tx_pin[216];
  assign mb1_FA1_TB0_IO_059_mb1_FB1_TB2_IO_073 = tx_pin[217];
  assign mb1_FA1_TB0_IO_060_mb1_FB1_TB2_IO_070 = tx_pin[218];
  assign mb1_FA1_TB0_IO_061_mb1_FB1_TB2_IO_071 = tx_pin[219];
  assign mb1_FA1_TB0_IO_062_mb1_FB1_TB2_IO_048 = tx_pin[220];
  assign mb1_FA1_TB0_IO_063_mb1_FB1_TB2_IO_049 = tx_pin[221];
  assign mb1_FA1_TB0_IO_064_mb1_FB1_TB2_IO_066 = tx_pin[222];
  assign mb1_FA1_TB0_IO_065_mb1_FB1_TB2_IO_067 = tx_pin[223];
  assign mb1_FA1_TB0_IO_066_mb1_FB1_TB2_IO_064 = tx_pin[224];
  assign mb1_FA1_TB0_IO_067_mb1_FB1_TB2_IO_065 = tx_pin[225];
  assign mb1_FA1_TB0_IO_068_mb1_FB1_TB2_IO_082 = tx_pin[226];
  assign mb1_FA1_TB0_IO_069_mb1_FB1_TB2_IO_083 = tx_pin[227];
  assign mb1_FA1_TB0_IO_070_mb1_FB1_TB2_IO_060 = tx_pin[228];
  assign mb1_FA1_TB0_IO_071_mb1_FB1_TB2_IO_061 = tx_pin[229];
  assign mb1_FA1_TB0_IO_072_mb1_FB1_TB2_IO_058 = tx_pin[230];
  assign mb1_FA1_TB0_IO_073_mb1_FB1_TB2_IO_059 = tx_pin[231];
  assign mb1_FA1_TB0_IO_074_mb1_FB1_TB2_IO_076 = tx_pin[232];
  assign mb1_FA1_TB0_IO_075_mb1_FB1_TB2_IO_077 = tx_pin[233];
  assign mb1_FA1_TB0_IO_076_mb1_FB1_TB2_IO_074 = tx_pin[234];
  assign mb1_FA1_TB0_IO_077_mb1_FB1_TB2_IO_075 = tx_pin[235];
  assign mb1_FA1_TB0_IO_078_mb1_FB1_TB2_IO_092 = tx_pin[236];
  assign mb1_FA1_TB0_IO_079_mb1_FB1_TB2_IO_093 = tx_pin[237];
  assign mb1_FA1_TB0_IO_080_mb1_FB1_TB2_IO_090 = tx_pin[238];
  assign mb1_FA1_TB0_IO_081_mb1_FB1_TB2_IO_091 = tx_pin[239];
  assign mb1_FA1_TB0_IO_082_mb1_FB1_TB2_IO_068 = tx_pin[240];
  assign mb1_FA1_TB0_IO_083_mb1_FB1_TB2_IO_069 = tx_pin[241];
  assign mb1_FA1_TB0_IO_084_mb1_FB1_TB2_IO_086 = tx_pin[242];
  assign mb1_FA1_TB0_IO_085_mb1_FB1_TB2_IO_087 = tx_pin[243];
  assign mb1_FA1_TB0_IO_086_mb1_FB1_TB2_IO_084 = tx_pin[244];
  assign mb1_FA1_TB0_IO_087_mb1_FB1_TB2_IO_085 = tx_pin[245];
  assign mb1_FA1_TB0_IO_088_mb1_FB1_TB2_IO_102 = tx_pin[246];
  assign mb1_FA1_TB0_IO_089_mb1_FB1_TB2_IO_103 = tx_pin[247];
  assign mb1_FA1_TB0_IO_090_mb1_FB1_TB2_IO_080 = tx_pin[248];
  assign mb1_FA1_TB0_IO_091_mb1_FB1_TB2_IO_081 = tx_pin[249];
  assign mb1_FA1_TB0_IO_092_mb1_FB1_TB2_IO_078 = tx_pin[250];
  assign mb1_FA1_TB0_IO_093_mb1_FB1_TB2_IO_079 = tx_pin[251];
  assign mb1_FA1_TB0_IO_094_mb1_FB1_TB2_IO_096 = tx_pin[252];
  assign mb1_FA1_TB0_IO_095_mb1_FB1_TB2_IO_097 = tx_pin[253];
  assign mb1_FA1_TB0_IO_096_mb1_FB1_TB2_IO_094 = tx_pin[254];
  assign mb1_FA1_TB0_IO_097_mb1_FB1_TB2_IO_095 = tx_pin[255];
  assign mb1_FA1_TB0_IO_098_mb1_FB1_TB2_IO_112 = tx_pin[256];
  assign mb1_FA1_TB0_IO_099_mb1_FB1_TB2_IO_113 = tx_pin[257];
  assign mb1_FA1_TB0_IO_100_mb1_FB1_TB2_IO_110 = tx_pin[258];
  assign mb1_FA1_TB0_IO_101_mb1_FB1_TB2_IO_111 = tx_pin[259];
  assign mb1_FA1_TB0_IO_102_mb1_FB1_TB2_IO_088 = tx_pin[260];
  assign mb1_FA1_TB0_IO_103_mb1_FB1_TB2_IO_089 = tx_pin[261];
  assign mb1_FA1_TB0_IO_104_mb1_FB1_TB2_IO_106 = tx_pin[262];
  assign mb1_FA1_TB0_IO_105_mb1_FB1_TB2_IO_107 = tx_pin[263];
  assign mb1_FA1_TB0_IO_106_mb1_FB1_TB2_IO_104 = tx_pin[264];
  assign mb1_FA1_TB0_IO_107_mb1_FB1_TB2_IO_105 = tx_pin[265];
  assign mb1_FA1_TB0_IO_108_mb1_FB1_TB2_IO_122 = tx_pin[266];
  assign mb1_FA1_TB0_IO_109_mb1_FB1_TB2_IO_123 = tx_pin[267];
  assign mb1_FA1_TB0_IO_110_mb1_FB1_TB2_IO_100 = tx_pin[268];
  assign mb1_FA1_TB0_IO_111_mb1_FB1_TB2_IO_101 = tx_pin[269];
  assign mb1_FA1_TB0_IO_112_mb1_FB1_TB2_IO_098 = tx_pin[270];
  assign mb1_FA1_TB0_IO_113_mb1_FB1_TB2_IO_099 = tx_pin[271];
  assign mb1_FA1_TB0_IO_114_mb1_FB1_TB2_IO_116 = tx_pin[272];
  assign mb1_FA1_TB0_IO_115_mb1_FB1_TB2_IO_117 = tx_pin[273];
  assign mb1_FA1_TB0_IO_116_mb1_FB1_TB2_IO_114 = tx_pin[274];
  assign mb1_FA1_TB0_IO_117_mb1_FB1_TB2_IO_115 = tx_pin[275];
  assign mb1_FA1_TB0_IO_118_mb1_FB1_TB2_IO_132 = tx_pin[276];
  assign mb1_FA1_TB0_IO_119_mb1_FB1_TB2_IO_133 = tx_pin[277];
  assign mb1_FA1_TB0_IO_120_mb1_FB1_TB2_IO_130 = tx_pin[278];
  assign mb1_FA1_TB0_IO_121_mb1_FB1_TB2_IO_131 = tx_pin[279];
  assign mb1_FA1_TB0_IO_122_mb1_FB1_TB2_IO_108 = tx_pin[280];
  assign mb1_FA1_TB0_IO_123_mb1_FB1_TB2_IO_109 = tx_pin[281];
  assign mb1_FA1_TB0_IO_124_mb1_FB1_TB2_IO_126 = tx_pin[282];
  assign mb1_FA1_TB0_IO_125_mb1_FB1_TB2_IO_127 = tx_pin[283];
  assign mb1_FA1_TB0_IO_126_mb1_FB1_TB2_IO_124 = tx_pin[284];
  assign mb1_FA1_TB0_IO_127_mb1_FB1_TB2_IO_125 = tx_pin[285];
  assign mb1_FA1_TB0_IO_130_mb1_FB1_TB2_IO_120 = tx_pin[286];
  assign mb1_FA1_TB0_IO_131_mb1_FB1_TB2_IO_121 = tx_pin[287];
  assign mb1_FA1_TB0_IO_132_mb1_FB1_TB2_IO_118 = tx_pin[288];
  assign mb1_FA1_TB0_IO_133_mb1_FB1_TB2_IO_119 = tx_pin[289];
  assign mb1_FA1_TB0_IO_134_mb1_FB1_TB2_IO_136 = tx_pin[290];
  assign mb1_FA1_TB0_IO_136_mb1_FB1_TB2_IO_134 = tx_pin[291];
  assign mb1_FA1_TB1_CLKIO_N_0_mb1_FB1_BB1_CLKIO_N_7 = tx_pin[292];
  assign mb1_FA1_TB1_CLKIO_N_1_mb1_FB1_BB1_CLKIO_N_6 = tx_pin[293];
  assign mb1_FA1_TB1_CLKIO_N_2_mb1_FB1_BB1_CLKIO_N_4 = tx_pin[294];
  assign mb1_FA1_TB1_CLKIO_N_3_mb1_FB1_BB1_CLKIO_N_3 = tx_pin[295];
  assign mb1_FA1_TB1_CLKIO_N_4_mb1_FB1_BB1_CLKIO_N_2 = tx_pin[296];
  assign mb1_FA1_TB1_CLKIO_N_5_mb1_FB1_BB1_IO_010 = tx_pin[297];
  assign mb1_FA1_TB1_CLKIO_N_6_mb1_FB1_BB1_CLKIO_N_1 = tx_pin[298];
  assign mb1_FA1_TB1_CLKIO_N_7_mb1_FB1_BB1_CLKIO_N_0 = tx_pin[299];
  assign mb1_FA1_TB1_CLKIO_P_0_mb1_FB1_BB1_CLKIO_P_7 = tx_pin[300];
  assign mb1_FA1_TB1_CLKIO_P_1_mb1_FB1_BB1_CLKIO_P_6 = tx_pin[301];
  assign mb1_FA1_TB1_CLKIO_P_2_mb1_FB1_BB1_CLKIO_P_4 = tx_pin[302];
  assign mb1_FA1_TB1_CLKIO_P_3_mb1_FB1_BB1_CLKIO_P_3 = tx_pin[303];
  assign mb1_FA1_TB1_CLKIO_P_4_mb1_FB1_BB1_CLKIO_P_2 = tx_pin[304];
  assign mb1_FA1_TB1_CLKIO_P_5_mb1_FB1_BB1_IO_011 = tx_pin[305];
  assign mb1_FA1_TB1_CLKIO_P_6_mb1_FB1_BB1_CLKIO_P_1 = tx_pin[306];
  assign mb1_FA1_TB1_CLKIO_P_7_mb1_FB1_BB1_CLKIO_P_0 = tx_pin[307];
  assign mb1_FA1_TB1_IO_004_mb1_FB1_BB1_IO_006 = tx_pin[308];
  assign mb1_FA1_TB1_IO_005_mb1_FB1_BB1_IO_007 = tx_pin[309];
  assign mb1_FA1_TB1_IO_006_mb1_FB1_BB1_IO_004 = tx_pin[310];
  assign mb1_FA1_TB1_IO_007_mb1_FB1_BB1_IO_005 = tx_pin[311];
  assign mb1_FA1_TB1_IO_008_mb1_FB1_BB1_IO_022 = tx_pin[312];
  assign mb1_FA1_TB1_IO_009_mb1_FB1_BB1_IO_023 = tx_pin[313];
  assign mb1_FA1_TB1_IO_010_mb1_FB1_BB1_CLKIO_N_5 = tx_pin[314];
  assign mb1_FA1_TB1_IO_011_mb1_FB1_BB1_CLKIO_P_5 = tx_pin[315];
  assign mb1_FA1_TB1_IO_012_mb1_FB1_BB1_IO_012 = tx_pin[316];
  assign mb1_FA1_TB1_IO_013_mb1_FB1_BB1_IO_013 = tx_pin[317];
  assign mb1_FA1_TB1_IO_014_mb1_FB1_BB1_IO_016 = tx_pin[318];
  assign mb1_FA1_TB1_IO_015_mb1_FB1_BB1_IO_017 = tx_pin[319];
  assign mb1_FA1_TB1_IO_016_mb1_FB1_BB1_IO_014 = tx_pin[320];
  assign mb1_FA1_TB1_IO_017_mb1_FB1_BB1_IO_015 = tx_pin[321];
  assign mb1_FA1_TB1_IO_018_mb1_FB1_BB1_IO_032 = tx_pin[322];
  assign mb1_FA1_TB1_IO_019_mb1_FB1_BB1_IO_033 = tx_pin[323];
  assign mb1_FA1_TB1_IO_020_mb1_FB1_BB1_IO_030 = tx_pin[324];
  assign mb1_FA1_TB1_IO_021_mb1_FB1_BB1_IO_031 = tx_pin[325];
  assign mb1_FA1_TB1_IO_022_mb1_FB1_BB1_IO_008 = tx_pin[326];
  assign mb1_FA1_TB1_IO_023_mb1_FB1_BB1_IO_009 = tx_pin[327];
  assign mb1_FA1_TB1_IO_024_mb1_FB1_BB1_IO_026 = tx_pin[328];
  assign mb1_FA1_TB1_IO_025_mb1_FB1_BB1_IO_027 = tx_pin[329];
  assign mb1_FA1_TB1_IO_026_mb1_FB1_BB1_IO_024 = tx_pin[330];
  assign mb1_FA1_TB1_IO_027_mb1_FB1_BB1_IO_025 = tx_pin[331];
  assign mb1_FA1_TB1_IO_028_mb1_FB1_BB1_IO_042 = tx_pin[332];
  assign mb1_FA1_TB1_IO_029_mb1_FB1_BB1_IO_043 = tx_pin[333];
  assign mb1_FA1_TB1_IO_030_mb1_FB1_BB1_IO_020 = tx_pin[334];
  assign mb1_FA1_TB1_IO_031_mb1_FB1_BB1_IO_021 = tx_pin[335];
  assign mb1_FA1_TB1_IO_032_mb1_FB1_BB1_IO_018 = tx_pin[336];
  assign mb1_FA1_TB1_IO_033_mb1_FB1_BB1_IO_019 = tx_pin[337];
  assign mb1_FA1_TB1_IO_034_mb1_FB1_BB1_IO_036 = tx_pin[338];
  assign mb1_FA1_TB1_IO_035_mb1_FB1_BB1_IO_037 = tx_pin[339];
  assign mb1_FA1_TB1_IO_036_mb1_FB1_BB1_IO_034 = tx_pin[340];
  assign mb1_FA1_TB1_IO_037_mb1_FB1_BB1_IO_035 = tx_pin[341];
  assign mb1_FA1_TB1_IO_038_mb1_FB1_BB1_IO_052 = tx_pin[342];
  assign mb1_FA1_TB1_IO_039_mb1_FB1_BB1_IO_053 = tx_pin[343];
  assign mb1_FA1_TB1_IO_040_mb1_FB1_BB1_IO_050 = tx_pin[344];
  assign mb1_FA1_TB1_IO_041_mb1_FB1_BB1_IO_051 = tx_pin[345];
  assign mb1_FA1_TB1_IO_042_mb1_FB1_BB1_IO_028 = tx_pin[346];
  assign mb1_FA1_TB1_IO_043_mb1_FB1_BB1_IO_029 = tx_pin[347];
  assign mb1_FA1_TB1_IO_044_mb1_FB1_BB1_IO_046 = tx_pin[348];
  assign mb1_FA1_TB1_IO_045_mb1_FB1_BB1_IO_047 = tx_pin[349];
  assign mb1_FA1_TB1_IO_046_mb1_FB1_BB1_IO_044 = tx_pin[350];
  assign mb1_FA1_TB1_IO_047_mb1_FB1_BB1_IO_045 = tx_pin[351];
  assign mb1_FA1_TB1_IO_048_mb1_FB1_BB1_IO_062 = tx_pin[352];
  assign mb1_FA1_TB1_IO_049_mb1_FB1_BB1_IO_063 = tx_pin[353];
  assign mb1_FA1_TB1_IO_050_mb1_FB1_BB1_IO_040 = tx_pin[354];
  assign mb1_FA1_TB1_IO_051_mb1_FB1_BB1_IO_041 = tx_pin[355];
  assign mb1_FA1_TB1_IO_052_mb1_FB1_BB1_IO_038 = tx_pin[356];
  assign mb1_FA1_TB1_IO_053_mb1_FB1_BB1_IO_039 = tx_pin[357];
  assign mb1_FA1_TB1_IO_054_mb1_FB1_BB1_IO_056 = tx_pin[358];
  assign mb1_FA1_TB1_IO_055_mb1_FB1_BB1_IO_057 = tx_pin[359];
  assign mb1_FA1_TB1_IO_056_mb1_FB1_BB1_IO_054 = tx_pin[360];
  assign mb1_FA1_TB1_IO_057_mb1_FB1_BB1_IO_055 = tx_pin[361];
  assign mb1_FA1_TB1_IO_058_mb1_FB1_BB1_IO_072 = tx_pin[362];
  assign mb1_FA1_TB1_IO_059_mb1_FB1_BB1_IO_073 = tx_pin[363];
  assign mb1_FA1_TB1_IO_060_mb1_FB1_BB1_IO_070 = tx_pin[364];
  assign mb1_FA1_TB1_IO_061_mb1_FB1_BB1_IO_071 = tx_pin[365];
  assign mb1_FA1_TB1_IO_062_mb1_FB1_BB1_IO_048 = tx_pin[366];
  assign mb1_FA1_TB1_IO_063_mb1_FB1_BB1_IO_049 = tx_pin[367];
  assign mb1_FA1_TB1_IO_064_mb1_FB1_BB1_IO_066 = tx_pin[368];
  assign mb1_FA1_TB1_IO_065_mb1_FB1_BB1_IO_067 = tx_pin[369];
  assign mb1_FA1_TB1_IO_066_mb1_FB1_BB1_IO_064 = tx_pin[370];
  assign mb1_FA1_TB1_IO_067_mb1_FB1_BB1_IO_065 = tx_pin[371];
  assign mb1_FA1_TB1_IO_068_mb1_FB1_BB1_IO_082 = tx_pin[372];
  assign mb1_FA1_TB1_IO_069_mb1_FB1_BB1_IO_083 = tx_pin[373];
  assign mb1_FA1_TB1_IO_070_mb1_FB1_BB1_IO_060 = tx_pin[374];
  assign mb1_FA1_TB1_IO_071_mb1_FB1_BB1_IO_061 = tx_pin[375];
  assign mb1_FA1_TB1_IO_072_mb1_FB1_BB1_IO_058 = tx_pin[376];
  assign mb1_FA1_TB1_IO_073_mb1_FB1_BB1_IO_059 = tx_pin[377];
  assign mb1_FA1_TB1_IO_074_mb1_FB1_BB1_IO_076 = tx_pin[378];
  assign mb1_FA1_TB1_IO_075_mb1_FB1_BB1_IO_077 = tx_pin[379];
  assign mb1_FA1_TB1_IO_076_mb1_FB1_BB1_IO_074 = tx_pin[380];
  assign mb1_FA1_TB1_IO_077_mb1_FB1_BB1_IO_075 = tx_pin[381];
  assign mb1_FA1_TB1_IO_078_mb1_FB1_BB1_IO_092 = tx_pin[382];
  assign mb1_FA1_TB1_IO_079_mb1_FB1_BB1_IO_093 = tx_pin[383];
  assign mb1_FA1_TB1_IO_080_mb1_FB1_BB1_IO_090 = tx_pin[384];
  assign mb1_FA1_TB1_IO_081_mb1_FB1_BB1_IO_091 = tx_pin[385];
  assign mb1_FA1_TB1_IO_082_mb1_FB1_BB1_IO_068 = tx_pin[386];
  assign mb1_FA1_TB1_IO_083_mb1_FB1_BB1_IO_069 = tx_pin[387];
  assign mb1_FA1_TB1_IO_084_mb1_FB1_BB1_IO_086 = tx_pin[388];
  assign mb1_FA1_TB1_IO_085_mb1_FB1_BB1_IO_087 = tx_pin[389];
  assign mb1_FA1_TB1_IO_086_mb1_FB1_BB1_IO_084 = tx_pin[390];
  assign mb1_FA1_TB1_IO_087_mb1_FB1_BB1_IO_085 = tx_pin[391];
  assign mb1_FA1_TB1_IO_088_mb1_FB1_BB1_IO_102 = tx_pin[392];
  assign mb1_FA1_TB1_IO_089_mb1_FB1_BB1_IO_103 = tx_pin[393];
  assign mb1_FA1_TB1_IO_090_mb1_FB1_BB1_IO_080 = tx_pin[394];
  assign mb1_FA1_TB1_IO_091_mb1_FB1_BB1_IO_081 = tx_pin[395];
  assign mb1_FA1_TB1_IO_092_mb1_FB1_BB1_IO_078 = tx_pin[396];
  assign mb1_FA1_TB1_IO_093_mb1_FB1_BB1_IO_079 = tx_pin[397];
  assign mb1_FA1_TB1_IO_094_mb1_FB1_BB1_IO_096 = tx_pin[398];
  assign mb1_FA1_TB1_IO_095_mb1_FB1_BB1_IO_097 = tx_pin[399];
  assign mb1_FA1_TB1_IO_096_mb1_FB1_BB1_IO_094 = tx_pin[400];
  assign mb1_FA1_TB1_IO_097_mb1_FB1_BB1_IO_095 = tx_pin[401];
  assign mb1_FA1_TB1_IO_098_mb1_FB1_BB1_IO_112 = tx_pin[402];
  assign mb1_FA1_TB1_IO_099_mb1_FB1_BB1_IO_113 = tx_pin[403];
  assign mb1_FA1_TB1_IO_100_mb1_FB1_BB1_IO_110 = tx_pin[404];
  assign mb1_FA1_TB1_IO_101_mb1_FB1_BB1_IO_111 = tx_pin[405];
  assign mb1_FA1_TB1_IO_102_mb1_FB1_BB1_IO_088 = tx_pin[406];
  assign mb1_FA1_TB1_IO_103_mb1_FB1_BB1_IO_089 = tx_pin[407];
  assign mb1_FA1_TB1_IO_104_mb1_FB1_BB1_IO_106 = tx_pin[408];
  assign mb1_FA1_TB1_IO_105_mb1_FB1_BB1_IO_107 = tx_pin[409];
  assign mb1_FA1_TB1_IO_106_mb1_FB1_BB1_IO_104 = tx_pin[410];
  assign mb1_FA1_TB1_IO_107_mb1_FB1_BB1_IO_105 = tx_pin[411];
  assign mb1_FA1_TB1_IO_108_mb1_FB1_BB1_IO_122 = tx_pin[412];
  assign mb1_FA1_TB1_IO_109_mb1_FB1_BB1_IO_123 = tx_pin[413];
  assign mb1_FA1_TB1_IO_110_mb1_FB1_BB1_IO_100 = tx_pin[414];
  assign mb1_FA1_TB1_IO_111_mb1_FB1_BB1_IO_101 = tx_pin[415];
  assign mb1_FA1_TB1_IO_112_mb1_FB1_BB1_IO_098 = tx_pin[416];
  assign mb1_FA1_TB1_IO_113_mb1_FB1_BB1_IO_099 = tx_pin[417];
  assign mb1_FA1_TB1_IO_114_mb1_FB1_BB1_IO_116 = tx_pin[418];
  assign mb1_FA1_TB1_IO_115_mb1_FB1_BB1_IO_117 = tx_pin[419];
  assign mb1_FA1_TB1_IO_116_mb1_FB1_BB1_IO_114 = tx_pin[420];
  assign mb1_FA1_TB1_IO_117_mb1_FB1_BB1_IO_115 = tx_pin[421];
  assign mb1_FA1_TB1_IO_118_mb1_FB1_BB1_IO_132 = tx_pin[422];
  assign mb1_FA1_TB1_IO_119_mb1_FB1_BB1_IO_133 = tx_pin[423];
  assign mb1_FA1_TB1_IO_120_mb1_FB1_BB1_IO_130 = tx_pin[424];
  assign mb1_FA1_TB1_IO_121_mb1_FB1_BB1_IO_131 = tx_pin[425];
  assign mb1_FA1_TB1_IO_122_mb1_FB1_BB1_IO_108 = tx_pin[426];
  assign mb1_FA1_TB1_IO_123_mb1_FB1_BB1_IO_109 = tx_pin[427];
  assign mb1_FA1_TB1_IO_124_mb1_FB1_BB1_IO_126 = tx_pin[428];
  assign mb1_FA1_TB1_IO_125_mb1_FB1_BB1_IO_127 = tx_pin[429];
  assign mb1_FA1_TB1_IO_126_mb1_FB1_BB1_IO_124 = tx_pin[430];
  assign mb1_FA1_TB1_IO_127_mb1_FB1_BB1_IO_125 = tx_pin[431];
  assign mb1_FA1_TB1_IO_130_mb1_FB1_BB1_IO_120 = tx_pin[432];
  assign mb1_FA1_TB1_IO_131_mb1_FB1_BB1_IO_121 = tx_pin[433];
  assign mb1_FA1_TB1_IO_132_mb1_FB1_BB1_IO_118 = tx_pin[434];
  assign mb1_FA1_TB1_IO_133_mb1_FB1_BB1_IO_119 = tx_pin[435];
  assign mb1_FA1_TB1_IO_134_mb1_FB1_BB1_IO_136 = tx_pin[436];
  assign mb1_FA1_TB1_IO_136_mb1_FB1_BB1_IO_134 = tx_pin[437];
  assign mb1_FA1_TB2_CLKIO_N_0_mb1_FB2_BB1_CLKIO_N_7 = tx_pin[438];
  assign mb1_FA1_TB2_CLKIO_N_1_mb1_FB2_BB1_CLKIO_N_6 = tx_pin[439];
  assign mb1_FA1_TB2_CLKIO_N_2_mb1_FB2_BB1_CLKIO_N_4 = tx_pin[440];
  assign mb1_FA1_TB2_CLKIO_N_3_mb1_FB2_BB1_CLKIO_N_3 = tx_pin[441];
  assign mb1_FA1_TB2_CLKIO_N_4_mb1_FB2_BB1_CLKIO_N_2 = tx_pin[442];
  assign mb1_FA1_TB2_CLKIO_N_5_mb1_FB2_BB1_IO_010 = tx_pin[443];
  assign mb1_FA1_TB2_CLKIO_N_6_mb1_FB2_BB1_CLKIO_N_1 = tx_pin[444];
  assign mb1_FA1_TB2_CLKIO_N_7_mb1_FB2_BB1_CLKIO_N_0 = tx_pin[445];
  assign mb1_FA1_TB2_CLKIO_P_0_mb1_FB2_BB1_CLKIO_P_7 = tx_pin[446];
  assign mb1_FA1_TB2_CLKIO_P_1_mb1_FB2_BB1_CLKIO_P_6 = tx_pin[447];
  assign mb1_FA1_TB2_CLKIO_P_2_mb1_FB2_BB1_CLKIO_P_4 = tx_pin[448];
  assign mb1_FA1_TB2_CLKIO_P_3_mb1_FB2_BB1_CLKIO_P_3 = tx_pin[449];
  assign mb1_FA1_TB2_CLKIO_P_4_mb1_FB2_BB1_CLKIO_P_2 = tx_pin[450];
  assign mb1_FA1_TB2_CLKIO_P_5_mb1_FB2_BB1_IO_011 = tx_pin[451];
  assign mb1_FA1_TB2_CLKIO_P_6_mb1_FB2_BB1_CLKIO_P_1 = tx_pin[452];
  assign mb1_FA1_TB2_CLKIO_P_7_mb1_FB2_BB1_CLKIO_P_0 = tx_pin[453];
  assign mb1_FA1_TB2_IO_004_mb1_FB2_BB1_IO_006 = tx_pin[454];
  assign mb1_FA1_TB2_IO_005_mb1_FB2_BB1_IO_007 = tx_pin[455];
  assign mb1_FA1_TB2_IO_006_mb1_FB2_BB1_IO_004 = tx_pin[456];
  assign mb1_FA1_TB2_IO_007_mb1_FB2_BB1_IO_005 = tx_pin[457];
  assign mb1_FA1_TB2_IO_008_mb1_FB2_BB1_IO_022 = tx_pin[458];
  assign mb1_FA1_TB2_IO_009_mb1_FB2_BB1_IO_023 = tx_pin[459];
  assign mb1_FA1_TB2_IO_010_mb1_FB2_BB1_CLKIO_N_5 = tx_pin[460];
  assign mb1_FA1_TB2_IO_011_mb1_FB2_BB1_CLKIO_P_5 = tx_pin[461];
  assign mb1_FA1_TB2_IO_012_mb1_FB2_BB1_IO_012 = tx_pin[462];
  assign mb1_FA1_TB2_IO_013_mb1_FB2_BB1_IO_013 = tx_pin[463];
  assign mb1_FA1_TB2_IO_014_mb1_FB2_BB1_IO_016 = tx_pin[464];
  assign mb1_FA1_TB2_IO_015_mb1_FB2_BB1_IO_017 = tx_pin[465];
  assign mb1_FA1_TB2_IO_016_mb1_FB2_BB1_IO_014 = tx_pin[466];
  assign mb1_FA1_TB2_IO_017_mb1_FB2_BB1_IO_015 = tx_pin[467];
  assign mb1_FA1_TB2_IO_018_mb1_FB2_BB1_IO_032 = tx_pin[468];
  assign mb1_FA1_TB2_IO_019_mb1_FB2_BB1_IO_033 = tx_pin[469];
  assign mb1_FA1_TB2_IO_020_mb1_FB2_BB1_IO_030 = tx_pin[470];
  assign mb1_FA1_TB2_IO_021_mb1_FB2_BB1_IO_031 = tx_pin[471];
  assign mb1_FA1_TB2_IO_022_mb1_FB2_BB1_IO_008 = tx_pin[472];
  assign mb1_FA1_TB2_IO_023_mb1_FB2_BB1_IO_009 = tx_pin[473];
  assign mb1_FA1_TB2_IO_024_mb1_FB2_BB1_IO_026 = tx_pin[474];
  assign mb1_FA1_TB2_IO_025_mb1_FB2_BB1_IO_027 = tx_pin[475];
  assign mb1_FA1_TB2_IO_026_mb1_FB2_BB1_IO_024 = tx_pin[476];
  assign mb1_FA1_TB2_IO_027_mb1_FB2_BB1_IO_025 = tx_pin[477];
  assign mb1_FA1_TB2_IO_028_mb1_FB2_BB1_IO_042 = tx_pin[478];
  assign mb1_FA1_TB2_IO_029_mb1_FB2_BB1_IO_043 = tx_pin[479];
  assign mb1_FA1_TB2_IO_030_mb1_FB2_BB1_IO_020 = tx_pin[480];
  assign mb1_FA1_TB2_IO_031_mb1_FB2_BB1_IO_021 = tx_pin[481];
  assign mb1_FA1_TB2_IO_032_mb1_FB2_BB1_IO_018 = tx_pin[482];
  assign mb1_FA1_TB2_IO_033_mb1_FB2_BB1_IO_019 = tx_pin[483];
  assign mb1_FA1_TB2_IO_034_mb1_FB2_BB1_IO_036 = tx_pin[484];
  assign mb1_FA1_TB2_IO_035_mb1_FB2_BB1_IO_037 = tx_pin[485];
  assign mb1_FA1_TB2_IO_036_mb1_FB2_BB1_IO_034 = tx_pin[486];
  assign mb1_FA1_TB2_IO_037_mb1_FB2_BB1_IO_035 = tx_pin[487];
  assign mb1_FA1_TB2_IO_038_mb1_FB2_BB1_IO_052 = tx_pin[488];
  assign mb1_FA1_TB2_IO_039_mb1_FB2_BB1_IO_053 = tx_pin[489];
  assign mb1_FA1_TB2_IO_040_mb1_FB2_BB1_IO_050 = tx_pin[490];
  assign mb1_FA1_TB2_IO_041_mb1_FB2_BB1_IO_051 = tx_pin[491];
  assign mb1_FA1_TB2_IO_042_mb1_FB2_BB1_IO_028 = tx_pin[492];
  assign mb1_FA1_TB2_IO_043_mb1_FB2_BB1_IO_029 = tx_pin[493];
  assign mb1_FA1_TB2_IO_044_mb1_FB2_BB1_IO_046 = tx_pin[494];
  assign mb1_FA1_TB2_IO_045_mb1_FB2_BB1_IO_047 = tx_pin[495];
  assign mb1_FA1_TB2_IO_046_mb1_FB2_BB1_IO_044 = tx_pin[496];
  assign mb1_FA1_TB2_IO_047_mb1_FB2_BB1_IO_045 = tx_pin[497];
  assign mb1_FA1_TB2_IO_048_mb1_FB2_BB1_IO_062 = tx_pin[498];
  assign mb1_FA1_TB2_IO_049_mb1_FB2_BB1_IO_063 = tx_pin[499];
  assign mb1_FA1_TB2_IO_050_mb1_FB2_BB1_IO_040 = tx_pin[500];
  assign mb1_FA1_TB2_IO_051_mb1_FB2_BB1_IO_041 = tx_pin[501];
  assign mb1_FA1_TB2_IO_052_mb1_FB2_BB1_IO_038 = tx_pin[502];
  assign mb1_FA1_TB2_IO_053_mb1_FB2_BB1_IO_039 = tx_pin[503];
  assign mb1_FA1_TB2_IO_054_mb1_FB2_BB1_IO_056 = tx_pin[504];
  assign mb1_FA1_TB2_IO_055_mb1_FB2_BB1_IO_057 = tx_pin[505];
  assign mb1_FA1_TB2_IO_056_mb1_FB2_BB1_IO_054 = tx_pin[506];
  assign mb1_FA1_TB2_IO_057_mb1_FB2_BB1_IO_055 = tx_pin[507];
  assign mb1_FA1_TB2_IO_058_mb1_FB2_BB1_IO_072 = tx_pin[508];
  assign mb1_FA1_TB2_IO_059_mb1_FB2_BB1_IO_073 = tx_pin[509];
  assign mb1_FA1_TB2_IO_060_mb1_FB2_BB1_IO_070 = tx_pin[510];
  assign mb1_FA1_TB2_IO_061_mb1_FB2_BB1_IO_071 = tx_pin[511];
  assign mb1_FA1_TB2_IO_062_mb1_FB2_BB1_IO_048 = tx_pin[512];
  assign mb1_FA1_TB2_IO_063_mb1_FB2_BB1_IO_049 = tx_pin[513];
  assign mb1_FA1_TB2_IO_064_mb1_FB2_BB1_IO_066 = tx_pin[514];
  assign mb1_FA1_TB2_IO_065_mb1_FB2_BB1_IO_067 = tx_pin[515];
  assign mb1_FA1_TB2_IO_066_mb1_FB2_BB1_IO_064 = tx_pin[516];
  assign mb1_FA1_TB2_IO_067_mb1_FB2_BB1_IO_065 = tx_pin[517];
  assign mb1_FA1_TB2_IO_068_mb1_FB2_BB1_IO_082 = tx_pin[518];
  assign mb1_FA1_TB2_IO_069_mb1_FB2_BB1_IO_083 = tx_pin[519];
  assign mb1_FA1_TB2_IO_070_mb1_FB2_BB1_IO_060 = tx_pin[520];
  assign mb1_FA1_TB2_IO_071_mb1_FB2_BB1_IO_061 = tx_pin[521];
  assign mb1_FA1_TB2_IO_072_mb1_FB2_BB1_IO_058 = tx_pin[522];
  assign mb1_FA1_TB2_IO_073_mb1_FB2_BB1_IO_059 = tx_pin[523];
  assign mb1_FA1_TB2_IO_074_mb1_FB2_BB1_IO_076 = tx_pin[524];
  assign mb1_FA1_TB2_IO_075_mb1_FB2_BB1_IO_077 = tx_pin[525];
  assign mb1_FA1_TB2_IO_076_mb1_FB2_BB1_IO_074 = tx_pin[526];
  assign mb1_FA1_TB2_IO_077_mb1_FB2_BB1_IO_075 = tx_pin[527];
  assign mb1_FA1_TB2_IO_078_mb1_FB2_BB1_IO_092 = tx_pin[528];
  assign mb1_FA1_TB2_IO_079_mb1_FB2_BB1_IO_093 = tx_pin[529];
  assign mb1_FA1_TB2_IO_080_mb1_FB2_BB1_IO_090 = tx_pin[530];
  assign mb1_FA1_TB2_IO_081_mb1_FB2_BB1_IO_091 = tx_pin[531];
  assign mb1_FA1_TB2_IO_082_mb1_FB2_BB1_IO_068 = tx_pin[532];
  assign mb1_FA1_TB2_IO_083_mb1_FB2_BB1_IO_069 = tx_pin[533];
  assign mb1_FA1_TB2_IO_084_mb1_FB2_BB1_IO_086 = tx_pin[534];
  assign mb1_FA1_TB2_IO_085_mb1_FB2_BB1_IO_087 = tx_pin[535];
  assign mb1_FA1_TB2_IO_086_mb1_FB2_BB1_IO_084 = tx_pin[536];
  assign mb1_FA1_TB2_IO_087_mb1_FB2_BB1_IO_085 = tx_pin[537];
  assign mb1_FA1_TB2_IO_088_mb1_FB2_BB1_IO_102 = tx_pin[538];
  assign mb1_FA1_TB2_IO_089_mb1_FB2_BB1_IO_103 = tx_pin[539];
  assign mb1_FA1_TB2_IO_090_mb1_FB2_BB1_IO_080 = tx_pin[540];
  assign mb1_FA1_TB2_IO_091_mb1_FB2_BB1_IO_081 = tx_pin[541];
  assign mb1_FA1_TB2_IO_092_mb1_FB2_BB1_IO_078 = tx_pin[542];
  assign mb1_FA1_TB2_IO_093_mb1_FB2_BB1_IO_079 = tx_pin[543];
  assign mb1_FA1_TB2_IO_094_mb1_FB2_BB1_IO_096 = tx_pin[544];
  assign mb1_FA1_TB2_IO_095_mb1_FB2_BB1_IO_097 = tx_pin[545];
  assign mb1_FA1_TB2_IO_096_mb1_FB2_BB1_IO_094 = tx_pin[546];
  assign mb1_FA1_TB2_IO_097_mb1_FB2_BB1_IO_095 = tx_pin[547];
  assign mb1_FA1_TB2_IO_098_mb1_FB2_BB1_IO_112 = tx_pin[548];
  assign mb1_FA1_TB2_IO_099_mb1_FB2_BB1_IO_113 = tx_pin[549];
  assign mb1_FA1_TB2_IO_100_mb1_FB2_BB1_IO_110 = tx_pin[550];
  assign mb1_FA1_TB2_IO_101_mb1_FB2_BB1_IO_111 = tx_pin[551];
  assign mb1_FA1_TB2_IO_102_mb1_FB2_BB1_IO_088 = tx_pin[552];
  assign mb1_FA1_TB2_IO_103_mb1_FB2_BB1_IO_089 = tx_pin[553];
  assign mb1_FA1_TB2_IO_104_mb1_FB2_BB1_IO_106 = tx_pin[554];
  assign mb1_FA1_TB2_IO_105_mb1_FB2_BB1_IO_107 = tx_pin[555];
  assign mb1_FA1_TB2_IO_106_mb1_FB2_BB1_IO_104 = tx_pin[556];
  assign mb1_FA1_TB2_IO_107_mb1_FB2_BB1_IO_105 = tx_pin[557];
  assign mb1_FA1_TB2_IO_108_mb1_FB2_BB1_IO_122 = tx_pin[558];
  assign mb1_FA1_TB2_IO_109_mb1_FB2_BB1_IO_123 = tx_pin[559];
  assign mb1_FA1_TB2_IO_110_mb1_FB2_BB1_IO_100 = tx_pin[560];
  assign mb1_FA1_TB2_IO_111_mb1_FB2_BB1_IO_101 = tx_pin[561];
  assign mb1_FA1_TB2_IO_112_mb1_FB2_BB1_IO_098 = tx_pin[562];
  assign mb1_FA1_TB2_IO_113_mb1_FB2_BB1_IO_099 = tx_pin[563];
  assign mb1_FA1_TB2_IO_114_mb1_FB2_BB1_IO_116 = tx_pin[564];
  assign mb1_FA1_TB2_IO_115_mb1_FB2_BB1_IO_117 = tx_pin[565];
  assign mb1_FA1_TB2_IO_116_mb1_FB2_BB1_IO_114 = tx_pin[566];
  assign mb1_FA1_TB2_IO_117_mb1_FB2_BB1_IO_115 = tx_pin[567];
  assign mb1_FA1_TB2_IO_118_mb1_FB2_BB1_IO_132 = tx_pin[568];
  assign mb1_FA1_TB2_IO_119_mb1_FB2_BB1_IO_133 = tx_pin[569];
  assign mb1_FA1_TB2_IO_120_mb1_FB2_BB1_IO_130 = tx_pin[570];
  assign mb1_FA1_TB2_IO_121_mb1_FB2_BB1_IO_131 = tx_pin[571];
  assign mb1_FA1_TB2_IO_122_mb1_FB2_BB1_IO_108 = tx_pin[572];
  assign mb1_FA1_TB2_IO_123_mb1_FB2_BB1_IO_109 = tx_pin[573];
  assign mb1_FA1_TB2_IO_124_mb1_FB2_BB1_IO_126 = tx_pin[574];
  assign mb1_FA1_TB2_IO_125_mb1_FB2_BB1_IO_127 = tx_pin[575];
  assign mb1_FA1_TB2_IO_126_mb1_FB2_BB1_IO_124 = tx_pin[576];
  assign mb1_FA1_TB2_IO_127_mb1_FB2_BB1_IO_125 = tx_pin[577];
  assign mb1_FA1_TB2_IO_130_mb1_FB2_BB1_IO_120 = tx_pin[578];
  assign mb1_FA1_TB2_IO_131_mb1_FB2_BB1_IO_121 = tx_pin[579];
  assign mb1_FA1_TB2_IO_132_mb1_FB2_BB1_IO_118 = tx_pin[580];
  assign mb1_FA1_TB2_IO_133_mb1_FB2_BB1_IO_119 = tx_pin[581];
  assign mb1_FA1_TB2_IO_134_mb1_FB2_BB1_IO_136 = tx_pin[582];
  assign mb1_FA1_TB2_IO_136_mb1_FB2_BB1_IO_134 = tx_pin[583];
  assign mb1_FA1_BA0_CLKIO_N_0_mb1_FB1_BA2_CLKIO_N_7 = tx_pin[584];
  assign mb1_FA1_BA0_CLKIO_N_1_mb1_FB1_BA2_CLKIO_N_6 = tx_pin[585];
  assign mb1_FA1_BA0_CLKIO_N_2_mb1_FB1_BA2_CLKIO_N_4 = tx_pin[586];
  assign mb1_FA1_BA0_CLKIO_N_3_mb1_FB1_BA2_CLKIO_N_3 = tx_pin[587];
  assign mb1_FA1_BA0_CLKIO_N_4_mb1_FB1_BA2_CLKIO_N_2 = tx_pin[588];
  assign mb1_FA1_BA0_CLKIO_N_5_mb1_FB1_BA2_IO_010 = tx_pin[589];
  assign mb1_FA1_BA0_CLKIO_N_6_mb1_FB1_BA2_CLKIO_N_1 = tx_pin[590];
  assign mb1_FA1_BA0_CLKIO_N_7_mb1_FB1_BA2_CLKIO_N_0 = tx_pin[591];
  assign mb1_FA1_BA0_CLKIO_P_0_mb1_FB1_BA2_CLKIO_P_7 = tx_pin[592];
  assign mb1_FA1_BA0_CLKIO_P_1_mb1_FB1_BA2_CLKIO_P_6 = tx_pin[593];
  assign mb1_FA1_BA0_CLKIO_P_2_mb1_FB1_BA2_CLKIO_P_4 = tx_pin[594];
  assign mb1_FA1_BA0_CLKIO_P_3_mb1_FB1_BA2_CLKIO_P_3 = tx_pin[595];
  assign mb1_FA1_BA0_CLKIO_P_4_mb1_FB1_BA2_CLKIO_P_2 = tx_pin[596];
  assign mb1_FA1_BA0_CLKIO_P_5_mb1_FB1_BA2_IO_011 = tx_pin[597];
  assign mb1_FA1_BA0_CLKIO_P_6_mb1_FB1_BA2_CLKIO_P_1 = tx_pin[598];
  assign mb1_FA1_BA0_CLKIO_P_7_mb1_FB1_BA2_CLKIO_P_0 = tx_pin[599];
  assign mb1_FA1_BA0_IO_004_mb1_FB1_BA2_IO_006 = tx_pin[600];
  assign mb1_FA1_BA0_IO_005_mb1_FB1_BA2_IO_007 = tx_pin[601];
  assign mb1_FA1_BA0_IO_006_mb1_FB1_BA2_IO_004 = tx_pin[602];
  assign mb1_FA1_BA0_IO_007_mb1_FB1_BA2_IO_005 = tx_pin[603];
  assign mb1_FA1_BA0_IO_008_mb1_FB1_BA2_IO_022 = tx_pin[604];
  assign mb1_FA1_BA0_IO_009_mb1_FB1_BA2_IO_023 = tx_pin[605];
  assign mb1_FA1_BA0_IO_010_mb1_FB1_BA2_CLKIO_N_5 = tx_pin[606];
  assign mb1_FA1_BA0_IO_011_mb1_FB1_BA2_CLKIO_P_5 = tx_pin[607];
  assign mb1_FA1_BA0_IO_012_mb1_FB1_BA2_IO_012 = tx_pin[608];
  assign mb1_FA1_BA0_IO_013_mb1_FB1_BA2_IO_013 = tx_pin[609];
  assign mb1_FA1_BA0_IO_014_mb1_FB1_BA2_IO_016 = tx_pin[610];
  assign mb1_FA1_BA0_IO_015_mb1_FB1_BA2_IO_017 = tx_pin[611];
  assign mb1_FA1_BA0_IO_016_mb1_FB1_BA2_IO_014 = tx_pin[612];
  assign mb1_FA1_BA0_IO_017_mb1_FB1_BA2_IO_015 = tx_pin[613];
  assign mb1_FA1_BA0_IO_018_mb1_FB1_BA2_IO_032 = tx_pin[614];
  assign mb1_FA1_BA0_IO_019_mb1_FB1_BA2_IO_033 = tx_pin[615];
  assign mb1_FA1_BA0_IO_020_mb1_FB1_BA2_IO_030 = tx_pin[616];
  assign mb1_FA1_BA0_IO_021_mb1_FB1_BA2_IO_031 = tx_pin[617];
  assign mb1_FA1_BA0_IO_022_mb1_FB1_BA2_IO_008 = tx_pin[618];
  assign mb1_FA1_BA0_IO_023_mb1_FB1_BA2_IO_009 = tx_pin[619];
  assign mb1_FA1_BA0_IO_024_mb1_FB1_BA2_IO_026 = tx_pin[620];
  assign mb1_FA1_BA0_IO_025_mb1_FB1_BA2_IO_027 = tx_pin[621];
  assign mb1_FA1_BA0_IO_026_mb1_FB1_BA2_IO_024 = tx_pin[622];
  assign mb1_FA1_BA0_IO_027_mb1_FB1_BA2_IO_025 = tx_pin[623];
  assign mb1_FA1_BA0_IO_028_mb1_FB1_BA2_IO_042 = tx_pin[624];
  assign mb1_FA1_BA0_IO_029_mb1_FB1_BA2_IO_043 = tx_pin[625];
  assign mb1_FA1_BA0_IO_030_mb1_FB1_BA2_IO_020 = tx_pin[626];
  assign mb1_FA1_BA0_IO_031_mb1_FB1_BA2_IO_021 = tx_pin[627];
  assign mb1_FA1_BA0_IO_032_mb1_FB1_BA2_IO_018 = tx_pin[628];
  assign mb1_FA1_BA0_IO_033_mb1_FB1_BA2_IO_019 = tx_pin[629];
  assign mb1_FA1_BA0_IO_034_mb1_FB1_BA2_IO_036 = tx_pin[630];
  assign mb1_FA1_BA0_IO_035_mb1_FB1_BA2_IO_037 = tx_pin[631];
  assign mb1_FA1_BA0_IO_036_mb1_FB1_BA2_IO_034 = tx_pin[632];
  assign mb1_FA1_BA0_IO_037_mb1_FB1_BA2_IO_035 = tx_pin[633];
  assign mb1_FA1_BA0_IO_038_mb1_FB1_BA2_IO_052 = tx_pin[634];
  assign mb1_FA1_BA0_IO_039_mb1_FB1_BA2_IO_053 = tx_pin[635];
  assign mb1_FA1_BA0_IO_040_mb1_FB1_BA2_IO_050 = tx_pin[636];
  assign mb1_FA1_BA0_IO_041_mb1_FB1_BA2_IO_051 = tx_pin[637];
  assign mb1_FA1_BA0_IO_042_mb1_FB1_BA2_IO_028 = tx_pin[638];
  assign mb1_FA1_BA0_IO_043_mb1_FB1_BA2_IO_029 = tx_pin[639];
  assign mb1_FA1_BA0_IO_044_mb1_FB1_BA2_IO_046 = tx_pin[640];
  assign mb1_FA1_BA0_IO_045_mb1_FB1_BA2_IO_047 = tx_pin[641];
  assign mb1_FA1_BA0_IO_046_mb1_FB1_BA2_IO_044 = tx_pin[642];
  assign mb1_FA1_BA0_IO_047_mb1_FB1_BA2_IO_045 = tx_pin[643];
  assign mb1_FA1_BA0_IO_048_mb1_FB1_BA2_IO_062 = tx_pin[644];
  assign mb1_FA1_BA0_IO_049_mb1_FB1_BA2_IO_063 = tx_pin[645];
  assign mb1_FA1_BA0_IO_050_mb1_FB1_BA2_IO_040 = tx_pin[646];
  assign mb1_FA1_BA0_IO_051_mb1_FB1_BA2_IO_041 = tx_pin[647];
  assign mb1_FA1_BA0_IO_052_mb1_FB1_BA2_IO_038 = tx_pin[648];
  assign mb1_FA1_BA0_IO_053_mb1_FB1_BA2_IO_039 = tx_pin[649];
  assign mb1_FA1_BA0_IO_054_mb1_FB1_BA2_IO_056 = tx_pin[650];
  assign mb1_FA1_BA0_IO_055_mb1_FB1_BA2_IO_057 = tx_pin[651];
  assign mb1_FA1_BA0_IO_056_mb1_FB1_BA2_IO_054 = tx_pin[652];
  assign mb1_FA1_BA0_IO_057_mb1_FB1_BA2_IO_055 = tx_pin[653];
  assign mb1_FA1_BA0_IO_058_mb1_FB1_BA2_IO_072 = tx_pin[654];
  assign mb1_FA1_BA0_IO_059_mb1_FB1_BA2_IO_073 = tx_pin[655];
  assign mb1_FA1_BA0_IO_060_mb1_FB1_BA2_IO_070 = tx_pin[656];
  assign mb1_FA1_BA0_IO_061_mb1_FB1_BA2_IO_071 = tx_pin[657];
  assign mb1_FA1_BA0_IO_062_mb1_FB1_BA2_IO_048 = tx_pin[658];
  assign mb1_FA1_BA0_IO_063_mb1_FB1_BA2_IO_049 = tx_pin[659];
  assign mb1_FA1_BA0_IO_064_mb1_FB1_BA2_IO_066 = tx_pin[660];
  assign mb1_FA1_BA0_IO_065_mb1_FB1_BA2_IO_067 = tx_pin[661];
  assign mb1_FA1_BA0_IO_066_mb1_FB1_BA2_IO_064 = tx_pin[662];
  assign mb1_FA1_BA0_IO_067_mb1_FB1_BA2_IO_065 = tx_pin[663];
  assign mb1_FA1_BA0_IO_068_mb1_FB1_BA2_IO_082 = tx_pin[664];
  assign mb1_FA1_BA0_IO_069_mb1_FB1_BA2_IO_083 = tx_pin[665];
  assign mb1_FA1_BA0_IO_070_mb1_FB1_BA2_IO_060 = tx_pin[666];
  assign mb1_FA1_BA0_IO_071_mb1_FB1_BA2_IO_061 = tx_pin[667];
  assign mb1_FA1_BA0_IO_072_mb1_FB1_BA2_IO_058 = tx_pin[668];
  assign mb1_FA1_BA0_IO_073_mb1_FB1_BA2_IO_059 = tx_pin[669];
  assign mb1_FA1_BA0_IO_074_mb1_FB1_BA2_IO_076 = tx_pin[670];
  assign mb1_FA1_BA0_IO_075_mb1_FB1_BA2_IO_077 = tx_pin[671];
  assign mb1_FA1_BA0_IO_076_mb1_FB1_BA2_IO_074 = tx_pin[672];
  assign mb1_FA1_BA0_IO_077_mb1_FB1_BA2_IO_075 = tx_pin[673];
  assign mb1_FA1_BA0_IO_078_mb1_FB1_BA2_IO_092 = tx_pin[674];
  assign mb1_FA1_BA0_IO_079_mb1_FB1_BA2_IO_093 = tx_pin[675];
  assign mb1_FA1_BA0_IO_080_mb1_FB1_BA2_IO_090 = tx_pin[676];
  assign mb1_FA1_BA0_IO_081_mb1_FB1_BA2_IO_091 = tx_pin[677];
  assign mb1_FA1_BA0_IO_082_mb1_FB1_BA2_IO_068 = tx_pin[678];
  assign mb1_FA1_BA0_IO_083_mb1_FB1_BA2_IO_069 = tx_pin[679];
  assign mb1_FA1_BA0_IO_084_mb1_FB1_BA2_IO_086 = tx_pin[680];
  assign mb1_FA1_BA0_IO_085_mb1_FB1_BA2_IO_087 = tx_pin[681];
  assign mb1_FA1_BA0_IO_086_mb1_FB1_BA2_IO_084 = tx_pin[682];
  assign mb1_FA1_BA0_IO_087_mb1_FB1_BA2_IO_085 = tx_pin[683];
  assign mb1_FA1_BA0_IO_088_mb1_FB1_BA2_IO_102 = tx_pin[684];
  assign mb1_FA1_BA0_IO_089_mb1_FB1_BA2_IO_103 = tx_pin[685];
  assign mb1_FA1_BA0_IO_090_mb1_FB1_BA2_IO_080 = tx_pin[686];
  assign mb1_FA1_BA0_IO_091_mb1_FB1_BA2_IO_081 = tx_pin[687];
  assign mb1_FA1_BA0_IO_092_mb1_FB1_BA2_IO_078 = tx_pin[688];
  assign mb1_FA1_BA0_IO_093_mb1_FB1_BA2_IO_079 = tx_pin[689];
  assign mb1_FA1_BA0_IO_094_mb1_FB1_BA2_IO_096 = tx_pin[690];
  assign mb1_FA1_BA0_IO_095_mb1_FB1_BA2_IO_097 = tx_pin[691];
  assign mb1_FA1_BA0_IO_096_mb1_FB1_BA2_IO_094 = tx_pin[692];
  assign mb1_FA1_BA0_IO_097_mb1_FB1_BA2_IO_095 = tx_pin[693];
  assign mb1_FA1_BA0_IO_098_mb1_FB1_BA2_IO_112 = tx_pin[694];
  assign mb1_FA1_BA0_IO_099_mb1_FB1_BA2_IO_113 = tx_pin[695];
  assign mb1_FA1_BA0_IO_100_mb1_FB1_BA2_IO_110 = tx_pin[696];
  assign mb1_FA1_BA0_IO_101_mb1_FB1_BA2_IO_111 = tx_pin[697];
  assign mb1_FA1_BA0_IO_102_mb1_FB1_BA2_IO_088 = tx_pin[698];
  assign mb1_FA1_BA0_IO_103_mb1_FB1_BA2_IO_089 = tx_pin[699];
  assign mb1_FA1_BA0_IO_104_mb1_FB1_BA2_IO_106 = tx_pin[700];
  assign mb1_FA1_BA0_IO_105_mb1_FB1_BA2_IO_107 = tx_pin[701];
  assign mb1_FA1_BA0_IO_106_mb1_FB1_BA2_IO_104 = tx_pin[702];
  assign mb1_FA1_BA0_IO_107_mb1_FB1_BA2_IO_105 = tx_pin[703];
  assign mb1_FA1_BA0_IO_108_mb1_FB1_BA2_IO_122 = tx_pin[704];
  assign mb1_FA1_BA0_IO_109_mb1_FB1_BA2_IO_123 = tx_pin[705];
  assign mb1_FA1_BA0_IO_110_mb1_FB1_BA2_IO_100 = tx_pin[706];
  assign mb1_FA1_BA0_IO_111_mb1_FB1_BA2_IO_101 = tx_pin[707];
  assign mb1_FA1_BA0_IO_112_mb1_FB1_BA2_IO_098 = tx_pin[708];
  assign mb1_FA1_BA0_IO_113_mb1_FB1_BA2_IO_099 = tx_pin[709];
  assign mb1_FA1_BA0_IO_114_mb1_FB1_BA2_IO_116 = tx_pin[710];
  assign mb1_FA1_BA0_IO_115_mb1_FB1_BA2_IO_117 = tx_pin[711];
  assign mb1_FA1_BA0_IO_116_mb1_FB1_BA2_IO_114 = tx_pin[712];
  assign mb1_FA1_BA0_IO_117_mb1_FB1_BA2_IO_115 = tx_pin[713];
  assign mb1_FA1_BA0_IO_118_mb1_FB1_BA2_IO_132 = tx_pin[714];
  assign mb1_FA1_BA0_IO_119_mb1_FB1_BA2_IO_133 = tx_pin[715];
  assign mb1_FA1_BA0_IO_120_mb1_FB1_BA2_IO_130 = tx_pin[716];
  assign mb1_FA1_BA0_IO_121_mb1_FB1_BA2_IO_131 = tx_pin[717];
  assign mb1_FA1_BA0_IO_122_mb1_FB1_BA2_IO_108 = tx_pin[718];
  assign mb1_FA1_BA0_IO_123_mb1_FB1_BA2_IO_109 = tx_pin[719];
  assign mb1_FA1_BA0_IO_124_mb1_FB1_BA2_IO_126 = tx_pin[720];
  assign mb1_FA1_BA0_IO_125_mb1_FB1_BA2_IO_127 = tx_pin[721];
  assign mb1_FA1_BA0_IO_126_mb1_FB1_BA2_IO_124 = tx_pin[722];
  assign mb1_FA1_BA0_IO_127_mb1_FB1_BA2_IO_125 = tx_pin[723];
  assign mb1_FA1_BA0_IO_130_mb1_FB1_BA2_IO_120 = tx_pin[724];
  assign mb1_FA1_BA0_IO_131_mb1_FB1_BA2_IO_121 = tx_pin[725];
  assign mb1_FA1_BA0_IO_132_mb1_FB1_BA2_IO_118 = tx_pin[726];
  assign mb1_FA1_BA0_IO_133_mb1_FB1_BA2_IO_119 = tx_pin[727];
  assign mb1_FA1_BA0_IO_134_mb1_FB1_BA2_IO_136 = tx_pin[728];
  assign mb1_FA1_BA0_IO_136_mb1_FB1_BA2_IO_134 = tx_pin[729];
  assign mb1_FA1_BA1_CLKIO_N_0_mb1_FA2_BB2_CLKIO_N_7 = tx_pin[730];
  assign mb1_FA1_BA1_CLKIO_N_1_mb1_FA2_BB2_CLKIO_N_6 = tx_pin[731];
  assign mb1_FA1_BA1_CLKIO_N_2_mb1_FA2_BB2_CLKIO_N_4 = tx_pin[732];
  assign mb1_FA1_BA1_CLKIO_N_3_mb1_FA2_BB2_CLKIO_N_3 = tx_pin[733];
  assign mb1_FA1_BA1_CLKIO_N_4_mb1_FA2_BB2_CLKIO_N_2 = tx_pin[734];
  assign mb1_FA1_BA1_CLKIO_N_5_mb1_FA2_BB2_IO_010 = tx_pin[735];
  assign mb1_FA1_BA1_CLKIO_N_6_mb1_FA2_BB2_CLKIO_N_1 = tx_pin[736];
  assign mb1_FA1_BA1_CLKIO_N_7_mb1_FA2_BB2_CLKIO_N_0 = tx_pin[737];
  assign mb1_FA1_BA1_CLKIO_P_0_mb1_FA2_BB2_CLKIO_P_7 = tx_pin[738];
  assign mb1_FA1_BA1_CLKIO_P_1_mb1_FA2_BB2_CLKIO_P_6 = tx_pin[739];
  assign mb1_FA1_BA1_CLKIO_P_2_mb1_FA2_BB2_CLKIO_P_4 = tx_pin[740];
  assign mb1_FA1_BA1_CLKIO_P_3_mb1_FA2_BB2_CLKIO_P_3 = tx_pin[741];
  assign mb1_FA1_BA1_CLKIO_P_4_mb1_FA2_BB2_CLKIO_P_2 = tx_pin[742];
  assign mb1_FA1_BA1_CLKIO_P_5_mb1_FA2_BB2_IO_011 = tx_pin[743];
  assign mb1_FA1_BA1_CLKIO_P_6_mb1_FA2_BB2_CLKIO_P_1 = tx_pin[744];
  assign mb1_FA1_BA1_CLKIO_P_7_mb1_FA2_BB2_CLKIO_P_0 = tx_pin[745];
  assign mb1_FA1_BA1_IO_004_mb1_FA2_BB2_IO_006 = tx_pin[746];
  assign mb1_FA1_BA1_IO_005_mb1_FA2_BB2_IO_007 = tx_pin[747];
  assign mb1_FA1_BA1_IO_006_mb1_FA2_BB2_IO_004 = tx_pin[748];
  assign mb1_FA1_BA1_IO_007_mb1_FA2_BB2_IO_005 = tx_pin[749];
  assign mb1_FA1_BA1_IO_008_mb1_FA2_BB2_IO_022 = tx_pin[750];
  assign mb1_FA1_BA1_IO_009_mb1_FA2_BB2_IO_023 = tx_pin[751];
  assign mb1_FA1_BA1_IO_010_mb1_FA2_BB2_CLKIO_N_5 = tx_pin[752];
  assign mb1_FA1_BA1_IO_011_mb1_FA2_BB2_CLKIO_P_5 = tx_pin[753];
  assign mb1_FA1_BA1_IO_012_mb1_FA2_BB2_IO_012 = tx_pin[754];
  assign mb1_FA1_BA1_IO_013_mb1_FA2_BB2_IO_013 = tx_pin[755];
  assign mb1_FA1_BA1_IO_014_mb1_FA2_BB2_IO_016 = tx_pin[756];
  assign mb1_FA1_BA1_IO_015_mb1_FA2_BB2_IO_017 = tx_pin[757];
  assign mb1_FA1_BA1_IO_016_mb1_FA2_BB2_IO_014 = tx_pin[758];
  assign mb1_FA1_BA1_IO_017_mb1_FA2_BB2_IO_015 = tx_pin[759];
  assign mb1_FA1_BA1_IO_018_mb1_FA2_BB2_IO_032 = tx_pin[760];
  assign mb1_FA1_BA1_IO_019_mb1_FA2_BB2_IO_033 = tx_pin[761];
  assign mb1_FA1_BA1_IO_020_mb1_FA2_BB2_IO_030 = tx_pin[762];
  assign mb1_FA1_BA1_IO_021_mb1_FA2_BB2_IO_031 = tx_pin[763];
  assign mb1_FA1_BA1_IO_022_mb1_FA2_BB2_IO_008 = tx_pin[764];
  assign mb1_FA1_BA1_IO_023_mb1_FA2_BB2_IO_009 = tx_pin[765];
  assign mb1_FA1_BA1_IO_024_mb1_FA2_BB2_IO_026 = tx_pin[766];
  assign mb1_FA1_BA1_IO_025_mb1_FA2_BB2_IO_027 = tx_pin[767];
  assign mb1_FA1_BA1_IO_026_mb1_FA2_BB2_IO_024 = tx_pin[768];
  assign mb1_FA1_BA1_IO_027_mb1_FA2_BB2_IO_025 = tx_pin[769];
  assign mb1_FA1_BA1_IO_028_mb1_FA2_BB2_IO_042 = tx_pin[770];
  assign mb1_FA1_BA1_IO_029_mb1_FA2_BB2_IO_043 = tx_pin[771];
  assign mb1_FA1_BA1_IO_030_mb1_FA2_BB2_IO_020 = tx_pin[772];
  assign mb1_FA1_BA1_IO_031_mb1_FA2_BB2_IO_021 = tx_pin[773];
  assign mb1_FA1_BA1_IO_032_mb1_FA2_BB2_IO_018 = tx_pin[774];
  assign mb1_FA1_BA1_IO_033_mb1_FA2_BB2_IO_019 = tx_pin[775];
  assign mb1_FA1_BA1_IO_034_mb1_FA2_BB2_IO_036 = tx_pin[776];
  assign mb1_FA1_BA1_IO_035_mb1_FA2_BB2_IO_037 = tx_pin[777];
  assign mb1_FA1_BA1_IO_036_mb1_FA2_BB2_IO_034 = tx_pin[778];
  assign mb1_FA1_BA1_IO_037_mb1_FA2_BB2_IO_035 = tx_pin[779];
  assign mb1_FA1_BA1_IO_038_mb1_FA2_BB2_IO_052 = tx_pin[780];
  assign mb1_FA1_BA1_IO_039_mb1_FA2_BB2_IO_053 = tx_pin[781];
  assign mb1_FA1_BA1_IO_040_mb1_FA2_BB2_IO_050 = tx_pin[782];
  assign mb1_FA1_BA1_IO_041_mb1_FA2_BB2_IO_051 = tx_pin[783];
  assign mb1_FA1_BA1_IO_042_mb1_FA2_BB2_IO_028 = tx_pin[784];
  assign mb1_FA1_BA1_IO_043_mb1_FA2_BB2_IO_029 = tx_pin[785];
  assign mb1_FA1_BA1_IO_044_mb1_FA2_BB2_IO_046 = tx_pin[786];
  assign mb1_FA1_BA1_IO_045_mb1_FA2_BB2_IO_047 = tx_pin[787];
  assign mb1_FA1_BA1_IO_046_mb1_FA2_BB2_IO_044 = tx_pin[788];
  assign mb1_FA1_BA1_IO_047_mb1_FA2_BB2_IO_045 = tx_pin[789];
  assign mb1_FA1_BA1_IO_048_mb1_FA2_BB2_IO_062 = tx_pin[790];
  assign mb1_FA1_BA1_IO_049_mb1_FA2_BB2_IO_063 = tx_pin[791];
  assign mb1_FA1_BA1_IO_050_mb1_FA2_BB2_IO_040 = tx_pin[792];
  assign mb1_FA1_BA1_IO_051_mb1_FA2_BB2_IO_041 = tx_pin[793];
  assign mb1_FA1_BA1_IO_052_mb1_FA2_BB2_IO_038 = tx_pin[794];
  assign mb1_FA1_BA1_IO_053_mb1_FA2_BB2_IO_039 = tx_pin[795];
  assign mb1_FA1_BA1_IO_054_mb1_FA2_BB2_IO_056 = tx_pin[796];
  assign mb1_FA1_BA1_IO_055_mb1_FA2_BB2_IO_057 = tx_pin[797];
  assign mb1_FA1_BA1_IO_056_mb1_FA2_BB2_IO_054 = tx_pin[798];
  assign mb1_FA1_BA1_IO_057_mb1_FA2_BB2_IO_055 = tx_pin[799];
  assign mb1_FA1_BA1_IO_058_mb1_FA2_BB2_IO_072 = tx_pin[800];
  assign mb1_FA1_BA1_IO_059_mb1_FA2_BB2_IO_073 = tx_pin[801];
  assign mb1_FA1_BA1_IO_060_mb1_FA2_BB2_IO_070 = tx_pin[802];
  assign mb1_FA1_BA1_IO_061_mb1_FA2_BB2_IO_071 = tx_pin[803];
  assign mb1_FA1_BA1_IO_062_mb1_FA2_BB2_IO_048 = tx_pin[804];
  assign mb1_FA1_BA1_IO_063_mb1_FA2_BB2_IO_049 = tx_pin[805];
  assign mb1_FA1_BA1_IO_064_mb1_FA2_BB2_IO_066 = tx_pin[806];
  assign mb1_FA1_BA1_IO_065_mb1_FA2_BB2_IO_067 = tx_pin[807];
  assign mb1_FA1_BA1_IO_066_mb1_FA2_BB2_IO_064 = tx_pin[808];
  assign mb1_FA1_BA1_IO_067_mb1_FA2_BB2_IO_065 = tx_pin[809];
  assign mb1_FA1_BA1_IO_068_mb1_FA2_BB2_IO_082 = tx_pin[810];
  assign mb1_FA1_BA1_IO_069_mb1_FA2_BB2_IO_083 = tx_pin[811];
  assign mb1_FA1_BA1_IO_070_mb1_FA2_BB2_IO_060 = tx_pin[812];
  assign mb1_FA1_BA1_IO_071_mb1_FA2_BB2_IO_061 = tx_pin[813];
  assign mb1_FA1_BA1_IO_072_mb1_FA2_BB2_IO_058 = tx_pin[814];
  assign mb1_FA1_BA1_IO_073_mb1_FA2_BB2_IO_059 = tx_pin[815];
  assign mb1_FA1_BA1_IO_074_mb1_FA2_BB2_IO_076 = tx_pin[816];
  assign mb1_FA1_BA1_IO_075_mb1_FA2_BB2_IO_077 = tx_pin[817];
  assign mb1_FA1_BA1_IO_076_mb1_FA2_BB2_IO_074 = tx_pin[818];
  assign mb1_FA1_BA1_IO_077_mb1_FA2_BB2_IO_075 = tx_pin[819];
  assign mb1_FA1_BA1_IO_078_mb1_FA2_BB2_IO_092 = tx_pin[820];
  assign mb1_FA1_BA1_IO_079_mb1_FA2_BB2_IO_093 = tx_pin[821];
  assign mb1_FA1_BA1_IO_080_mb1_FA2_BB2_IO_090 = tx_pin[822];
  assign mb1_FA1_BA1_IO_081_mb1_FA2_BB2_IO_091 = tx_pin[823];
  assign mb1_FA1_BA1_IO_082_mb1_FA2_BB2_IO_068 = tx_pin[824];
  assign mb1_FA1_BA1_IO_083_mb1_FA2_BB2_IO_069 = tx_pin[825];
  assign mb1_FA1_BA1_IO_084_mb1_FA2_BB2_IO_086 = tx_pin[826];
  assign mb1_FA1_BA1_IO_085_mb1_FA2_BB2_IO_087 = tx_pin[827];
  assign mb1_FA1_BA1_IO_086_mb1_FA2_BB2_IO_084 = tx_pin[828];
  assign mb1_FA1_BA1_IO_087_mb1_FA2_BB2_IO_085 = tx_pin[829];
  assign mb1_FA1_BA1_IO_088_mb1_FA2_BB2_IO_102 = tx_pin[830];
  assign mb1_FA1_BA1_IO_089_mb1_FA2_BB2_IO_103 = tx_pin[831];
  assign mb1_FA1_BA1_IO_090_mb1_FA2_BB2_IO_080 = tx_pin[832];
  assign mb1_FA1_BA1_IO_091_mb1_FA2_BB2_IO_081 = tx_pin[833];
  assign mb1_FA1_BA1_IO_092_mb1_FA2_BB2_IO_078 = tx_pin[834];
  assign mb1_FA1_BA1_IO_093_mb1_FA2_BB2_IO_079 = tx_pin[835];
  assign mb1_FA1_BA1_IO_094_mb1_FA2_BB2_IO_096 = tx_pin[836];
  assign mb1_FA1_BA1_IO_095_mb1_FA2_BB2_IO_097 = tx_pin[837];
  assign mb1_FA1_BA1_IO_096_mb1_FA2_BB2_IO_094 = tx_pin[838];
  assign mb1_FA1_BA1_IO_097_mb1_FA2_BB2_IO_095 = tx_pin[839];
  assign mb1_FA1_BA1_IO_098_mb1_FA2_BB2_IO_112 = tx_pin[840];
  assign mb1_FA1_BA1_IO_099_mb1_FA2_BB2_IO_113 = tx_pin[841];
  assign mb1_FA1_BA1_IO_100_mb1_FA2_BB2_IO_110 = tx_pin[842];
  assign mb1_FA1_BA1_IO_101_mb1_FA2_BB2_IO_111 = tx_pin[843];
  assign mb1_FA1_BA1_IO_102_mb1_FA2_BB2_IO_088 = tx_pin[844];
  assign mb1_FA1_BA1_IO_103_mb1_FA2_BB2_IO_089 = tx_pin[845];
  assign mb1_FA1_BA1_IO_104_mb1_FA2_BB2_IO_106 = tx_pin[846];
  assign mb1_FA1_BA1_IO_105_mb1_FA2_BB2_IO_107 = tx_pin[847];
  assign mb1_FA1_BA1_IO_106_mb1_FA2_BB2_IO_104 = tx_pin[848];
  assign mb1_FA1_BA1_IO_107_mb1_FA2_BB2_IO_105 = tx_pin[849];
  assign mb1_FA1_BA1_IO_108_mb1_FA2_BB2_IO_122 = tx_pin[850];
  assign mb1_FA1_BA1_IO_109_mb1_FA2_BB2_IO_123 = tx_pin[851];
  assign mb1_FA1_BA1_IO_110_mb1_FA2_BB2_IO_100 = tx_pin[852];
  assign mb1_FA1_BA1_IO_111_mb1_FA2_BB2_IO_101 = tx_pin[853];
  assign mb1_FA1_BA1_IO_112_mb1_FA2_BB2_IO_098 = tx_pin[854];
  assign mb1_FA1_BA1_IO_113_mb1_FA2_BB2_IO_099 = tx_pin[855];
  assign mb1_FA1_BA1_IO_114_mb1_FA2_BB2_IO_116 = tx_pin[856];
  assign mb1_FA1_BA1_IO_115_mb1_FA2_BB2_IO_117 = tx_pin[857];
  assign mb1_FA1_BA1_IO_116_mb1_FA2_BB2_IO_114 = tx_pin[858];
  assign mb1_FA1_BA1_IO_117_mb1_FA2_BB2_IO_115 = tx_pin[859];
  assign mb1_FA1_BA1_IO_118_mb1_FA2_BB2_IO_132 = tx_pin[860];
  assign mb1_FA1_BA1_IO_119_mb1_FA2_BB2_IO_133 = tx_pin[861];
  assign mb1_FA1_BA1_IO_120_mb1_FA2_BB2_IO_130 = tx_pin[862];
  assign mb1_FA1_BA1_IO_121_mb1_FA2_BB2_IO_131 = tx_pin[863];
  assign mb1_FA1_BA1_IO_122_mb1_FA2_BB2_IO_108 = tx_pin[864];
  assign mb1_FA1_BA1_IO_123_mb1_FA2_BB2_IO_109 = tx_pin[865];
  assign mb1_FA1_BA1_IO_124_mb1_FA2_BB2_IO_126 = tx_pin[866];
  assign mb1_FA1_BA1_IO_125_mb1_FA2_BB2_IO_127 = tx_pin[867];
  assign mb1_FA1_BA1_IO_126_mb1_FA2_BB2_IO_124 = tx_pin[868];
  assign mb1_FA1_BA1_IO_127_mb1_FA2_BB2_IO_125 = tx_pin[869];
  assign mb1_FA1_BA1_IO_130_mb1_FA2_BB2_IO_120 = tx_pin[870];
  assign mb1_FA1_BA1_IO_131_mb1_FA2_BB2_IO_121 = tx_pin[871];
  assign mb1_FA1_BA1_IO_132_mb1_FA2_BB2_IO_118 = tx_pin[872];
  assign mb1_FA1_BA1_IO_133_mb1_FA2_BB2_IO_119 = tx_pin[873];
  assign mb1_FA1_BA1_IO_134_mb1_FA2_BB2_IO_136 = tx_pin[874];
  assign mb1_FA1_BA1_IO_136_mb1_FA2_BB2_IO_134 = tx_pin[875];
  assign mb1_FA1_BA2_CLKIO_N_0_mb1_FB1_BB0_CLKIO_N_7 = tx_pin[876];
  assign mb1_FA1_BA2_CLKIO_N_1_mb1_FB1_BB0_CLKIO_N_6 = tx_pin[877];
  assign mb1_FA1_BA2_CLKIO_N_2_mb1_FB1_BB0_CLKIO_N_4 = tx_pin[878];
  assign mb1_FA1_BA2_CLKIO_N_3_mb1_FB1_BB0_CLKIO_N_3 = tx_pin[879];
  assign mb1_FA1_BA2_CLKIO_N_4_mb1_FB1_BB0_CLKIO_N_2 = tx_pin[880];
  assign mb1_FA1_BA2_CLKIO_N_5_mb1_FB1_BB0_IO_010 = tx_pin[881];
  assign mb1_FA1_BA2_CLKIO_N_6_mb1_FB1_BB0_CLKIO_N_1 = tx_pin[882];
  assign mb1_FA1_BA2_CLKIO_N_7_mb1_FB1_BB0_CLKIO_N_0 = tx_pin[883];
  assign mb1_FA1_BA2_CLKIO_P_0_mb1_FB1_BB0_CLKIO_P_7 = tx_pin[884];
  assign mb1_FA1_BA2_CLKIO_P_1_mb1_FB1_BB0_CLKIO_P_6 = tx_pin[885];
  assign mb1_FA1_BA2_CLKIO_P_2_mb1_FB1_BB0_CLKIO_P_4 = tx_pin[886];
  assign mb1_FA1_BA2_CLKIO_P_3_mb1_FB1_BB0_CLKIO_P_3 = tx_pin[887];
  assign mb1_FA1_BA2_CLKIO_P_4_mb1_FB1_BB0_CLKIO_P_2 = tx_pin[888];
  assign mb1_FA1_BA2_CLKIO_P_5_mb1_FB1_BB0_IO_011 = tx_pin[889];
  assign mb1_FA1_BA2_CLKIO_P_6_mb1_FB1_BB0_CLKIO_P_1 = tx_pin[890];
  assign mb1_FA1_BA2_CLKIO_P_7_mb1_FB1_BB0_CLKIO_P_0 = tx_pin[891];
  assign mb1_FA1_BA2_IO_004_mb1_FB1_BB0_IO_006 = tx_pin[892];
  assign mb1_FA1_BA2_IO_005_mb1_FB1_BB0_IO_007 = tx_pin[893];
  assign mb1_FA1_BA2_IO_006_mb1_FB1_BB0_IO_004 = tx_pin[894];
  assign mb1_FA1_BA2_IO_007_mb1_FB1_BB0_IO_005 = tx_pin[895];
  assign mb1_FA1_BA2_IO_008_mb1_FB1_BB0_IO_022 = tx_pin[896];
  assign mb1_FA1_BA2_IO_009_mb1_FB1_BB0_IO_023 = tx_pin[897];
  assign mb1_FA1_BA2_IO_010_mb1_FB1_BB0_CLKIO_N_5 = tx_pin[898];
  assign mb1_FA1_BA2_IO_011_mb1_FB1_BB0_CLKIO_P_5 = tx_pin[899];
  assign mb1_FA1_BA2_IO_012_mb1_FB1_BB0_IO_012 = tx_pin[900];
  assign mb1_FA1_BA2_IO_013_mb1_FB1_BB0_IO_013 = tx_pin[901];
  assign mb1_FA1_BA2_IO_014_mb1_FB1_BB0_IO_016 = tx_pin[902];
  assign mb1_FA1_BA2_IO_015_mb1_FB1_BB0_IO_017 = tx_pin[903];
  assign mb1_FA1_BA2_IO_016_mb1_FB1_BB0_IO_014 = tx_pin[904];
  assign mb1_FA1_BA2_IO_017_mb1_FB1_BB0_IO_015 = tx_pin[905];
  assign mb1_FA1_BA2_IO_018_mb1_FB1_BB0_IO_032 = tx_pin[906];
  assign mb1_FA1_BA2_IO_019_mb1_FB1_BB0_IO_033 = tx_pin[907];
  assign mb1_FA1_BA2_IO_020_mb1_FB1_BB0_IO_030 = tx_pin[908];
  assign mb1_FA1_BA2_IO_021_mb1_FB1_BB0_IO_031 = tx_pin[909];
  assign mb1_FA1_BA2_IO_022_mb1_FB1_BB0_IO_008 = tx_pin[910];
  assign mb1_FA1_BA2_IO_023_mb1_FB1_BB0_IO_009 = tx_pin[911];
  assign mb1_FA1_BA2_IO_024_mb1_FB1_BB0_IO_026 = tx_pin[912];
  assign mb1_FA1_BA2_IO_025_mb1_FB1_BB0_IO_027 = tx_pin[913];
  assign mb1_FA1_BA2_IO_026_mb1_FB1_BB0_IO_024 = tx_pin[914];
  assign mb1_FA1_BA2_IO_027_mb1_FB1_BB0_IO_025 = tx_pin[915];
  assign mb1_FA1_BA2_IO_028_mb1_FB1_BB0_IO_042 = tx_pin[916];
  assign mb1_FA1_BA2_IO_029_mb1_FB1_BB0_IO_043 = tx_pin[917];
  assign mb1_FA1_BA2_IO_030_mb1_FB1_BB0_IO_020 = tx_pin[918];
  assign mb1_FA1_BA2_IO_031_mb1_FB1_BB0_IO_021 = tx_pin[919];
  assign mb1_FA1_BA2_IO_032_mb1_FB1_BB0_IO_018 = tx_pin[920];
  assign mb1_FA1_BA2_IO_033_mb1_FB1_BB0_IO_019 = tx_pin[921];
  assign mb1_FA1_BA2_IO_034_mb1_FB1_BB0_IO_036 = tx_pin[922];
  assign mb1_FA1_BA2_IO_035_mb1_FB1_BB0_IO_037 = tx_pin[923];
  assign mb1_FA1_BA2_IO_036_mb1_FB1_BB0_IO_034 = tx_pin[924];
  assign mb1_FA1_BA2_IO_037_mb1_FB1_BB0_IO_035 = tx_pin[925];
  assign mb1_FA1_BA2_IO_038_mb1_FB1_BB0_IO_052 = tx_pin[926];
  assign mb1_FA1_BA2_IO_039_mb1_FB1_BB0_IO_053 = tx_pin[927];
  assign mb1_FA1_BA2_IO_040_mb1_FB1_BB0_IO_050 = tx_pin[928];
  assign mb1_FA1_BA2_IO_041_mb1_FB1_BB0_IO_051 = tx_pin[929];
  assign mb1_FA1_BA2_IO_042_mb1_FB1_BB0_IO_028 = tx_pin[930];
  assign mb1_FA1_BA2_IO_043_mb1_FB1_BB0_IO_029 = tx_pin[931];
  assign mb1_FA1_BA2_IO_044_mb1_FB1_BB0_IO_046 = tx_pin[932];
  assign mb1_FA1_BA2_IO_045_mb1_FB1_BB0_IO_047 = tx_pin[933];
  assign mb1_FA1_BA2_IO_046_mb1_FB1_BB0_IO_044 = tx_pin[934];
  assign mb1_FA1_BA2_IO_047_mb1_FB1_BB0_IO_045 = tx_pin[935];
  assign mb1_FA1_BA2_IO_048_mb1_FB1_BB0_IO_062 = tx_pin[936];
  assign mb1_FA1_BA2_IO_049_mb1_FB1_BB0_IO_063 = tx_pin[937];
  assign mb1_FA1_BA2_IO_050_mb1_FB1_BB0_IO_040 = tx_pin[938];
  assign mb1_FA1_BA2_IO_051_mb1_FB1_BB0_IO_041 = tx_pin[939];
  assign mb1_FA1_BA2_IO_052_mb1_FB1_BB0_IO_038 = tx_pin[940];
  assign mb1_FA1_BA2_IO_053_mb1_FB1_BB0_IO_039 = tx_pin[941];
  assign mb1_FA1_BA2_IO_054_mb1_FB1_BB0_IO_056 = tx_pin[942];
  assign mb1_FA1_BA2_IO_055_mb1_FB1_BB0_IO_057 = tx_pin[943];
  assign mb1_FA1_BA2_IO_056_mb1_FB1_BB0_IO_054 = tx_pin[944];
  assign mb1_FA1_BA2_IO_057_mb1_FB1_BB0_IO_055 = tx_pin[945];
  assign mb1_FA1_BA2_IO_058_mb1_FB1_BB0_IO_072 = tx_pin[946];
  assign mb1_FA1_BA2_IO_059_mb1_FB1_BB0_IO_073 = tx_pin[947];
  assign mb1_FA1_BA2_IO_060_mb1_FB1_BB0_IO_070 = tx_pin[948];
  assign mb1_FA1_BA2_IO_061_mb1_FB1_BB0_IO_071 = tx_pin[949];
  assign mb1_FA1_BA2_IO_062_mb1_FB1_BB0_IO_048 = tx_pin[950];
  assign mb1_FA1_BA2_IO_063_mb1_FB1_BB0_IO_049 = tx_pin[951];
  assign mb1_FA1_BA2_IO_064_mb1_FB1_BB0_IO_066 = tx_pin[952];
  assign mb1_FA1_BA2_IO_065_mb1_FB1_BB0_IO_067 = tx_pin[953];
  assign mb1_FA1_BA2_IO_066_mb1_FB1_BB0_IO_064 = tx_pin[954];
  assign mb1_FA1_BA2_IO_067_mb1_FB1_BB0_IO_065 = tx_pin[955];
  assign mb1_FA1_BA2_IO_068_mb1_FB1_BB0_IO_082 = tx_pin[956];
  assign mb1_FA1_BA2_IO_069_mb1_FB1_BB0_IO_083 = tx_pin[957];
  assign mb1_FA1_BA2_IO_070_mb1_FB1_BB0_IO_060 = tx_pin[958];
  assign mb1_FA1_BA2_IO_071_mb1_FB1_BB0_IO_061 = tx_pin[959];
  assign mb1_FA1_BA2_IO_072_mb1_FB1_BB0_IO_058 = tx_pin[960];
  assign mb1_FA1_BA2_IO_073_mb1_FB1_BB0_IO_059 = tx_pin[961];
  assign mb1_FA1_BA2_IO_074_mb1_FB1_BB0_IO_076 = tx_pin[962];
  assign mb1_FA1_BA2_IO_075_mb1_FB1_BB0_IO_077 = tx_pin[963];
  assign mb1_FA1_BA2_IO_076_mb1_FB1_BB0_IO_074 = tx_pin[964];
  assign mb1_FA1_BA2_IO_077_mb1_FB1_BB0_IO_075 = tx_pin[965];
  assign mb1_FA1_BA2_IO_078_mb1_FB1_BB0_IO_092 = tx_pin[966];
  assign mb1_FA1_BA2_IO_079_mb1_FB1_BB0_IO_093 = tx_pin[967];
  assign mb1_FA1_BA2_IO_080_mb1_FB1_BB0_IO_090 = tx_pin[968];
  assign mb1_FA1_BA2_IO_081_mb1_FB1_BB0_IO_091 = tx_pin[969];
  assign mb1_FA1_BA2_IO_082_mb1_FB1_BB0_IO_068 = tx_pin[970];
  assign mb1_FA1_BA2_IO_083_mb1_FB1_BB0_IO_069 = tx_pin[971];
  assign mb1_FA1_BA2_IO_084_mb1_FB1_BB0_IO_086 = tx_pin[972];
  assign mb1_FA1_BA2_IO_085_mb1_FB1_BB0_IO_087 = tx_pin[973];
  assign mb1_FA1_BA2_IO_086_mb1_FB1_BB0_IO_084 = tx_pin[974];
  assign mb1_FA1_BA2_IO_087_mb1_FB1_BB0_IO_085 = tx_pin[975];
  assign mb1_FA1_BA2_IO_088_mb1_FB1_BB0_IO_102 = tx_pin[976];
  assign mb1_FA1_BA2_IO_089_mb1_FB1_BB0_IO_103 = tx_pin[977];
  assign mb1_FA1_BA2_IO_090_mb1_FB1_BB0_IO_080 = tx_pin[978];
  assign mb1_FA1_BA2_IO_091_mb1_FB1_BB0_IO_081 = tx_pin[979];
  assign mb1_FA1_BA2_IO_092_mb1_FB1_BB0_IO_078 = tx_pin[980];
  assign mb1_FA1_BA2_IO_093_mb1_FB1_BB0_IO_079 = tx_pin[981];
  assign mb1_FA1_BA2_IO_094_mb1_FB1_BB0_IO_096 = tx_pin[982];
  assign mb1_FA1_BA2_IO_095_mb1_FB1_BB0_IO_097 = tx_pin[983];
  assign mb1_FA1_BA2_IO_096_mb1_FB1_BB0_IO_094 = tx_pin[984];
  assign mb1_FA1_BA2_IO_097_mb1_FB1_BB0_IO_095 = tx_pin[985];
  assign mb1_FA1_BA2_IO_098_mb1_FB1_BB0_IO_112 = tx_pin[986];
  assign mb1_FA1_BA2_IO_099_mb1_FB1_BB0_IO_113 = tx_pin[987];
  assign mb1_FA1_BA2_IO_100_mb1_FB1_BB0_IO_110 = tx_pin[988];
  assign mb1_FA1_BA2_IO_101_mb1_FB1_BB0_IO_111 = tx_pin[989];
  assign mb1_FA1_BA2_IO_102_mb1_FB1_BB0_IO_088 = tx_pin[990];
  assign mb1_FA1_BA2_IO_103_mb1_FB1_BB0_IO_089 = tx_pin[991];
  assign mb1_FA1_BA2_IO_104_mb1_FB1_BB0_IO_106 = tx_pin[992];
  assign mb1_FA1_BA2_IO_105_mb1_FB1_BB0_IO_107 = tx_pin[993];
  assign mb1_FA1_BA2_IO_106_mb1_FB1_BB0_IO_104 = tx_pin[994];
  assign mb1_FA1_BA2_IO_107_mb1_FB1_BB0_IO_105 = tx_pin[995];
  assign mb1_FA1_BA2_IO_108_mb1_FB1_BB0_IO_122 = tx_pin[996];
  assign mb1_FA1_BA2_IO_109_mb1_FB1_BB0_IO_123 = tx_pin[997];
  assign mb1_FA1_BA2_IO_110_mb1_FB1_BB0_IO_100 = tx_pin[998];
  assign mb1_FA1_BA2_IO_111_mb1_FB1_BB0_IO_101 = tx_pin[999];
  assign mb1_FA1_BA2_IO_112_mb1_FB1_BB0_IO_098 = tx_pin[1000];
  assign mb1_FA1_BA2_IO_113_mb1_FB1_BB0_IO_099 = tx_pin[1001];
  assign mb1_FA1_BA2_IO_114_mb1_FB1_BB0_IO_116 = tx_pin[1002];
  assign mb1_FA1_BA2_IO_115_mb1_FB1_BB0_IO_117 = tx_pin[1003];
  assign mb1_FA1_BA2_IO_116_mb1_FB1_BB0_IO_114 = tx_pin[1004];
  assign mb1_FA1_BA2_IO_117_mb1_FB1_BB0_IO_115 = tx_pin[1005];
  assign mb1_FA1_BA2_IO_118_mb1_FB1_BB0_IO_132 = tx_pin[1006];
  assign mb1_FA1_BA2_IO_119_mb1_FB1_BB0_IO_133 = tx_pin[1007];
  assign mb1_FA1_BA2_IO_120_mb1_FB1_BB0_IO_130 = tx_pin[1008];
  assign mb1_FA1_BA2_IO_121_mb1_FB1_BB0_IO_131 = tx_pin[1009];
  assign mb1_FA1_BA2_IO_122_mb1_FB1_BB0_IO_108 = tx_pin[1010];
  assign mb1_FA1_BA2_IO_123_mb1_FB1_BB0_IO_109 = tx_pin[1011];
  assign mb1_FA1_BA2_IO_124_mb1_FB1_BB0_IO_126 = tx_pin[1012];
  assign mb1_FA1_BA2_IO_125_mb1_FB1_BB0_IO_127 = tx_pin[1013];
  assign mb1_FA1_BA2_IO_126_mb1_FB1_BB0_IO_124 = tx_pin[1014];
  assign mb1_FA1_BA2_IO_127_mb1_FB1_BB0_IO_125 = tx_pin[1015];
  assign mb1_FA1_BA2_IO_130_mb1_FB1_BB0_IO_120 = tx_pin[1016];
  assign mb1_FA1_BA2_IO_131_mb1_FB1_BB0_IO_121 = tx_pin[1017];
  assign mb1_FA1_BA2_IO_132_mb1_FB1_BB0_IO_118 = tx_pin[1018];
  assign mb1_FA1_BA2_IO_133_mb1_FB1_BB0_IO_119 = tx_pin[1019];
  assign mb1_FA1_BA2_IO_134_mb1_FB1_BB0_IO_136 = tx_pin[1020];
  assign mb1_FA1_BA2_IO_136_mb1_FB1_BB0_IO_134 = tx_pin[1021];
  assign mb1_FA1_BB0_CLKIO_N_0_mb1_FB1_BB2_CLKIO_N_7 = tx_pin[1022];
  assign mb1_FA1_BB0_CLKIO_N_1_mb1_FB1_BB2_CLKIO_N_6 = tx_pin[1023];
  assign mb1_FA1_BB0_CLKIO_N_2_mb1_FB1_BB2_CLKIO_N_4 = tx_pin[1024];
  assign mb1_FA1_BB0_CLKIO_N_3_mb1_FB1_BB2_CLKIO_N_3 = tx_pin[1025];
  assign mb1_FA1_BB0_CLKIO_N_4_mb1_FB1_BB2_CLKIO_N_2 = tx_pin[1026];
  assign mb1_FA1_BB0_CLKIO_N_5_mb1_FB1_BB2_IO_010 = tx_pin[1027];
  assign mb1_FA1_BB0_CLKIO_N_6_mb1_FB1_BB2_CLKIO_N_1 = tx_pin[1028];
  assign mb1_FA1_BB0_CLKIO_N_7_mb1_FB1_BB2_CLKIO_N_0 = tx_pin[1029];
  assign mb1_FA1_BB0_CLKIO_P_0_mb1_FB1_BB2_CLKIO_P_7 = tx_pin[1030];
  assign mb1_FA1_BB0_CLKIO_P_1_mb1_FB1_BB2_CLKIO_P_6 = tx_pin[1031];
  assign mb1_FA1_BB0_CLKIO_P_2_mb1_FB1_BB2_CLKIO_P_4 = tx_pin[1032];
  assign mb1_FA1_BB0_CLKIO_P_3_mb1_FB1_BB2_CLKIO_P_3 = tx_pin[1033];
  assign mb1_FA1_BB0_CLKIO_P_4_mb1_FB1_BB2_CLKIO_P_2 = tx_pin[1034];
  assign mb1_FA1_BB0_CLKIO_P_5_mb1_FB1_BB2_IO_011 = tx_pin[1035];
  assign mb1_FA1_BB0_CLKIO_P_6_mb1_FB1_BB2_CLKIO_P_1 = tx_pin[1036];
  assign mb1_FA1_BB0_CLKIO_P_7_mb1_FB1_BB2_CLKIO_P_0 = tx_pin[1037];
  assign mb1_FA1_BB0_IO_004_mb1_FB1_BB2_IO_006 = tx_pin[1038];
  assign mb1_FA1_BB0_IO_005_mb1_FB1_BB2_IO_007 = tx_pin[1039];
  assign mb1_FA1_BB0_IO_006_mb1_FB1_BB2_IO_004 = tx_pin[1040];
  assign mb1_FA1_BB0_IO_007_mb1_FB1_BB2_IO_005 = tx_pin[1041];
  assign mb1_FA1_BB0_IO_008_mb1_FB1_BB2_IO_022 = tx_pin[1042];
  assign mb1_FA1_BB0_IO_009_mb1_FB1_BB2_IO_023 = tx_pin[1043];
  assign mb1_FA1_BB0_IO_010_mb1_FB1_BB2_CLKIO_N_5 = tx_pin[1044];
  assign mb1_FA1_BB0_IO_011_mb1_FB1_BB2_CLKIO_P_5 = tx_pin[1045];
  assign mb1_FA1_BB0_IO_012_mb1_FB1_BB2_IO_012 = tx_pin[1046];
  assign mb1_FA1_BB0_IO_013_mb1_FB1_BB2_IO_013 = tx_pin[1047];
  assign mb1_FA1_BB0_IO_014_mb1_FB1_BB2_IO_016 = tx_pin[1048];
  assign mb1_FA1_BB0_IO_015_mb1_FB1_BB2_IO_017 = tx_pin[1049];
  assign mb1_FA1_BB0_IO_016_mb1_FB1_BB2_IO_014 = tx_pin[1050];
  assign mb1_FA1_BB0_IO_017_mb1_FB1_BB2_IO_015 = tx_pin[1051];
  assign mb1_FA1_BB0_IO_018_mb1_FB1_BB2_IO_032 = tx_pin[1052];
  assign mb1_FA1_BB0_IO_019_mb1_FB1_BB2_IO_033 = tx_pin[1053];
  assign mb1_FA1_BB0_IO_020_mb1_FB1_BB2_IO_030 = tx_pin[1054];
  assign mb1_FA1_BB0_IO_021_mb1_FB1_BB2_IO_031 = tx_pin[1055];
  assign mb1_FA1_BB0_IO_022_mb1_FB1_BB2_IO_008 = tx_pin[1056];
  assign mb1_FA1_BB0_IO_023_mb1_FB1_BB2_IO_009 = tx_pin[1057];
  assign mb1_FA1_BB0_IO_024_mb1_FB1_BB2_IO_026 = tx_pin[1058];
  assign mb1_FA1_BB0_IO_025_mb1_FB1_BB2_IO_027 = tx_pin[1059];
  assign mb1_FA1_BB0_IO_026_mb1_FB1_BB2_IO_024 = tx_pin[1060];
  assign mb1_FA1_BB0_IO_027_mb1_FB1_BB2_IO_025 = tx_pin[1061];
  assign mb1_FA1_BB0_IO_028_mb1_FB1_BB2_IO_042 = tx_pin[1062];
  assign mb1_FA1_BB0_IO_029_mb1_FB1_BB2_IO_043 = tx_pin[1063];
  assign mb1_FA1_BB0_IO_030_mb1_FB1_BB2_IO_020 = tx_pin[1064];
  assign mb1_FA1_BB0_IO_031_mb1_FB1_BB2_IO_021 = tx_pin[1065];
  assign mb1_FA1_BB0_IO_032_mb1_FB1_BB2_IO_018 = tx_pin[1066];
  assign mb1_FA1_BB0_IO_033_mb1_FB1_BB2_IO_019 = tx_pin[1067];
  assign mb1_FA1_BB0_IO_034_mb1_FB1_BB2_IO_036 = tx_pin[1068];
  assign mb1_FA1_BB0_IO_035_mb1_FB1_BB2_IO_037 = tx_pin[1069];
  assign mb1_FA1_BB0_IO_036_mb1_FB1_BB2_IO_034 = tx_pin[1070];
  assign mb1_FA1_BB0_IO_037_mb1_FB1_BB2_IO_035 = tx_pin[1071];
  assign mb1_FA1_BB0_IO_038_mb1_FB1_BB2_IO_052 = tx_pin[1072];
  assign mb1_FA1_BB0_IO_039_mb1_FB1_BB2_IO_053 = tx_pin[1073];
  assign mb1_FA1_BB0_IO_040_mb1_FB1_BB2_IO_050 = tx_pin[1074];
  assign mb1_FA1_BB0_IO_041_mb1_FB1_BB2_IO_051 = tx_pin[1075];
  assign mb1_FA1_BB0_IO_042_mb1_FB1_BB2_IO_028 = tx_pin[1076];
  assign mb1_FA1_BB0_IO_043_mb1_FB1_BB2_IO_029 = tx_pin[1077];
  assign mb1_FA1_BB0_IO_044_mb1_FB1_BB2_IO_046 = tx_pin[1078];
  assign mb1_FA1_BB0_IO_045_mb1_FB1_BB2_IO_047 = tx_pin[1079];
  assign mb1_FA1_BB0_IO_046_mb1_FB1_BB2_IO_044 = tx_pin[1080];
  assign mb1_FA1_BB0_IO_047_mb1_FB1_BB2_IO_045 = tx_pin[1081];
  assign mb1_FA1_BB0_IO_048_mb1_FB1_BB2_IO_062 = tx_pin[1082];
  assign mb1_FA1_BB0_IO_049_mb1_FB1_BB2_IO_063 = tx_pin[1083];
  assign mb1_FA1_BB0_IO_050_mb1_FB1_BB2_IO_040 = tx_pin[1084];
  assign mb1_FA1_BB0_IO_051_mb1_FB1_BB2_IO_041 = tx_pin[1085];
  assign mb1_FA1_BB0_IO_052_mb1_FB1_BB2_IO_038 = tx_pin[1086];
  assign mb1_FA1_BB0_IO_053_mb1_FB1_BB2_IO_039 = tx_pin[1087];
  assign mb1_FA1_BB0_IO_054_mb1_FB1_BB2_IO_056 = tx_pin[1088];
  assign mb1_FA1_BB0_IO_055_mb1_FB1_BB2_IO_057 = tx_pin[1089];
  assign mb1_FA1_BB0_IO_056_mb1_FB1_BB2_IO_054 = tx_pin[1090];
  assign mb1_FA1_BB0_IO_057_mb1_FB1_BB2_IO_055 = tx_pin[1091];
  assign mb1_FA1_BB0_IO_058_mb1_FB1_BB2_IO_072 = tx_pin[1092];
  assign mb1_FA1_BB0_IO_059_mb1_FB1_BB2_IO_073 = tx_pin[1093];
  assign mb1_FA1_BB0_IO_060_mb1_FB1_BB2_IO_070 = tx_pin[1094];
  assign mb1_FA1_BB0_IO_061_mb1_FB1_BB2_IO_071 = tx_pin[1095];
  assign mb1_FA1_BB0_IO_062_mb1_FB1_BB2_IO_048 = tx_pin[1096];
  assign mb1_FA1_BB0_IO_063_mb1_FB1_BB2_IO_049 = tx_pin[1097];
  assign mb1_FA1_BB0_IO_064_mb1_FB1_BB2_IO_066 = tx_pin[1098];
  assign mb1_FA1_BB0_IO_065_mb1_FB1_BB2_IO_067 = tx_pin[1099];
  assign mb1_FA1_BB0_IO_066_mb1_FB1_BB2_IO_064 = tx_pin[1100];
  assign mb1_FA1_BB0_IO_067_mb1_FB1_BB2_IO_065 = tx_pin[1101];
  assign mb1_FA1_BB0_IO_068_mb1_FB1_BB2_IO_082 = tx_pin[1102];
  assign mb1_FA1_BB0_IO_069_mb1_FB1_BB2_IO_083 = tx_pin[1103];
  assign mb1_FA1_BB0_IO_070_mb1_FB1_BB2_IO_060 = tx_pin[1104];
  assign mb1_FA1_BB0_IO_071_mb1_FB1_BB2_IO_061 = tx_pin[1105];
  assign mb1_FA1_BB0_IO_072_mb1_FB1_BB2_IO_058 = tx_pin[1106];
  assign mb1_FA1_BB0_IO_073_mb1_FB1_BB2_IO_059 = tx_pin[1107];
  assign mb1_FA1_BB0_IO_074_mb1_FB1_BB2_IO_076 = tx_pin[1108];
  assign mb1_FA1_BB0_IO_075_mb1_FB1_BB2_IO_077 = tx_pin[1109];
  assign mb1_FA1_BB0_IO_076_mb1_FB1_BB2_IO_074 = tx_pin[1110];
  assign mb1_FA1_BB0_IO_077_mb1_FB1_BB2_IO_075 = tx_pin[1111];
  assign mb1_FA1_BB0_IO_078_mb1_FB1_BB2_IO_092 = tx_pin[1112];
  assign mb1_FA1_BB0_IO_079_mb1_FB1_BB2_IO_093 = tx_pin[1113];
  assign mb1_FA1_BB0_IO_080_mb1_FB1_BB2_IO_090 = tx_pin[1114];
  assign mb1_FA1_BB0_IO_081_mb1_FB1_BB2_IO_091 = tx_pin[1115];
  assign mb1_FA1_BB0_IO_082_mb1_FB1_BB2_IO_068 = tx_pin[1116];
  assign mb1_FA1_BB0_IO_083_mb1_FB1_BB2_IO_069 = tx_pin[1117];
  assign mb1_FA1_BB0_IO_084_mb1_FB1_BB2_IO_086 = tx_pin[1118];
  assign mb1_FA1_BB0_IO_085_mb1_FB1_BB2_IO_087 = tx_pin[1119];
  assign mb1_FA1_BB0_IO_086_mb1_FB1_BB2_IO_084 = tx_pin[1120];
  assign mb1_FA1_BB0_IO_087_mb1_FB1_BB2_IO_085 = tx_pin[1121];
  assign mb1_FA1_BB0_IO_088_mb1_FB1_BB2_IO_102 = tx_pin[1122];
  assign mb1_FA1_BB0_IO_089_mb1_FB1_BB2_IO_103 = tx_pin[1123];
  assign mb1_FA1_BB0_IO_090_mb1_FB1_BB2_IO_080 = tx_pin[1124];
  assign mb1_FA1_BB0_IO_091_mb1_FB1_BB2_IO_081 = tx_pin[1125];
  assign mb1_FA1_BB0_IO_092_mb1_FB1_BB2_IO_078 = tx_pin[1126];
  assign mb1_FA1_BB0_IO_093_mb1_FB1_BB2_IO_079 = tx_pin[1127];
  assign mb1_FA1_BB0_IO_094_mb1_FB1_BB2_IO_096 = tx_pin[1128];
  assign mb1_FA1_BB0_IO_095_mb1_FB1_BB2_IO_097 = tx_pin[1129];
  assign mb1_FA1_BB0_IO_096_mb1_FB1_BB2_IO_094 = tx_pin[1130];
  assign mb1_FA1_BB0_IO_097_mb1_FB1_BB2_IO_095 = tx_pin[1131];
  assign mb1_FA1_BB0_IO_098_mb1_FB1_BB2_IO_112 = tx_pin[1132];
  assign mb1_FA1_BB0_IO_099_mb1_FB1_BB2_IO_113 = tx_pin[1133];
  assign mb1_FA1_BB0_IO_100_mb1_FB1_BB2_IO_110 = tx_pin[1134];
  assign mb1_FA1_BB0_IO_101_mb1_FB1_BB2_IO_111 = tx_pin[1135];
  assign mb1_FA1_BB0_IO_102_mb1_FB1_BB2_IO_088 = tx_pin[1136];
  assign mb1_FA1_BB0_IO_103_mb1_FB1_BB2_IO_089 = tx_pin[1137];
  assign mb1_FA1_BB0_IO_104_mb1_FB1_BB2_IO_106 = tx_pin[1138];
  assign mb1_FA1_BB0_IO_105_mb1_FB1_BB2_IO_107 = tx_pin[1139];
  assign mb1_FA1_BB0_IO_106_mb1_FB1_BB2_IO_104 = tx_pin[1140];
  assign mb1_FA1_BB0_IO_107_mb1_FB1_BB2_IO_105 = tx_pin[1141];
  assign mb1_FA1_BB0_IO_108_mb1_FB1_BB2_IO_122 = tx_pin[1142];
  assign mb1_FA1_BB0_IO_109_mb1_FB1_BB2_IO_123 = tx_pin[1143];
  assign mb1_FA1_BB0_IO_110_mb1_FB1_BB2_IO_100 = tx_pin[1144];
  assign mb1_FA1_BB0_IO_111_mb1_FB1_BB2_IO_101 = tx_pin[1145];
  assign mb1_FA1_BB0_IO_112_mb1_FB1_BB2_IO_098 = tx_pin[1146];
  assign mb1_FA1_BB0_IO_113_mb1_FB1_BB2_IO_099 = tx_pin[1147];
  assign mb1_FA1_BB0_IO_114_mb1_FB1_BB2_IO_116 = tx_pin[1148];
  assign mb1_FA1_BB0_IO_115_mb1_FB1_BB2_IO_117 = tx_pin[1149];
  assign mb1_FA1_BB0_IO_116_mb1_FB1_BB2_IO_114 = tx_pin[1150];
  assign mb1_FA1_BB0_IO_117_mb1_FB1_BB2_IO_115 = tx_pin[1151];
  assign mb1_FA1_BB0_IO_118_mb1_FB1_BB2_IO_132 = tx_pin[1152];
  assign mb1_FA1_BB0_IO_119_mb1_FB1_BB2_IO_133 = tx_pin[1153];
  assign mb1_FA1_BB0_IO_120_mb1_FB1_BB2_IO_130 = tx_pin[1154];
  assign mb1_FA1_BB0_IO_121_mb1_FB1_BB2_IO_131 = tx_pin[1155];
  assign mb1_FA1_BB0_IO_122_mb1_FB1_BB2_IO_108 = tx_pin[1156];
  assign mb1_FA1_BB0_IO_123_mb1_FB1_BB2_IO_109 = tx_pin[1157];
  assign mb1_FA1_BB0_IO_124_mb1_FB1_BB2_IO_126 = tx_pin[1158];
  assign mb1_FA1_BB0_IO_125_mb1_FB1_BB2_IO_127 = tx_pin[1159];
  assign mb1_FA1_BB0_IO_126_mb1_FB1_BB2_IO_124 = tx_pin[1160];
  assign mb1_FA1_BB0_IO_127_mb1_FB1_BB2_IO_125 = tx_pin[1161];
  assign mb1_FA1_BB0_IO_130_mb1_FB1_BB2_IO_120 = tx_pin[1162];
  assign mb1_FA1_BB0_IO_131_mb1_FB1_BB2_IO_121 = tx_pin[1163];
  assign mb1_FA1_BB0_IO_132_mb1_FB1_BB2_IO_118 = tx_pin[1164];
  assign mb1_FA1_BB0_IO_133_mb1_FB1_BB2_IO_119 = tx_pin[1165];
  assign mb1_FA1_BB0_IO_134_mb1_FB1_BB2_IO_136 = tx_pin[1166];
  assign mb1_FA1_BB0_IO_136_mb1_FB1_BB2_IO_134 = tx_pin[1167];
  assign mb1_FA1_BB1_CLKIO_N_0_mb1_FA2_BB1_CLKIO_N_7 = tx_pin[1168];
  assign mb1_FA1_BB1_CLKIO_N_1_mb1_FA2_BB1_CLKIO_N_6 = tx_pin[1169];
  assign mb1_FA1_BB1_CLKIO_N_2_mb1_FA2_BB1_CLKIO_N_4 = tx_pin[1170];
  assign mb1_FA1_BB1_CLKIO_N_3_mb1_FA2_BB1_CLKIO_N_3 = tx_pin[1171];
  assign mb1_FA1_BB1_CLKIO_N_4_mb1_FA2_BB1_CLKIO_N_2 = tx_pin[1172];
  assign mb1_FA1_BB1_CLKIO_N_5_mb1_FA2_BB1_IO_010 = tx_pin[1173];
  assign mb1_FA1_BB1_CLKIO_N_6_mb1_FA2_BB1_CLKIO_N_1 = tx_pin[1174];
  assign mb1_FA1_BB1_CLKIO_N_7_mb1_FA2_BB1_CLKIO_N_0 = tx_pin[1175];
  assign mb1_FA1_BB1_CLKIO_P_0_mb1_FA2_BB1_CLKIO_P_7 = tx_pin[1176];
  assign mb1_FA1_BB1_CLKIO_P_1_mb1_FA2_BB1_CLKIO_P_6 = tx_pin[1177];
  assign mb1_FA1_BB1_CLKIO_P_2_mb1_FA2_BB1_CLKIO_P_4 = tx_pin[1178];
  assign mb1_FA1_BB1_CLKIO_P_3_mb1_FA2_BB1_CLKIO_P_3 = tx_pin[1179];
  assign mb1_FA1_BB1_CLKIO_P_4_mb1_FA2_BB1_CLKIO_P_2 = tx_pin[1180];
  assign mb1_FA1_BB1_CLKIO_P_5_mb1_FA2_BB1_IO_011 = tx_pin[1181];
  assign mb1_FA1_BB1_CLKIO_P_6_mb1_FA2_BB1_CLKIO_P_1 = tx_pin[1182];
  assign mb1_FA1_BB1_CLKIO_P_7_mb1_FA2_BB1_CLKIO_P_0 = tx_pin[1183];
  assign mb1_FA1_BB1_IO_004_mb1_FA2_BB1_IO_006 = tx_pin[1184];
  assign mb1_FA1_BB1_IO_005_mb1_FA2_BB1_IO_007 = tx_pin[1185];
  assign mb1_FA1_BB1_IO_006_mb1_FA2_BB1_IO_004 = tx_pin[1186];
  assign mb1_FA1_BB1_IO_007_mb1_FA2_BB1_IO_005 = tx_pin[1187];
  assign mb1_FA1_BB1_IO_008_mb1_FA2_BB1_IO_022 = tx_pin[1188];
  assign mb1_FA1_BB1_IO_009_mb1_FA2_BB1_IO_023 = tx_pin[1189];
  assign mb1_FA1_BB1_IO_010_mb1_FA2_BB1_CLKIO_N_5 = tx_pin[1190];
  assign mb1_FA1_BB1_IO_011_mb1_FA2_BB1_CLKIO_P_5 = tx_pin[1191];
  assign mb1_FA1_BB1_IO_012_mb1_FA2_BB1_IO_012 = tx_pin[1192];
  assign mb1_FA1_BB1_IO_013_mb1_FA2_BB1_IO_013 = tx_pin[1193];
  assign mb1_FA1_BB1_IO_014_mb1_FA2_BB1_IO_016 = tx_pin[1194];
  assign mb1_FA1_BB1_IO_015_mb1_FA2_BB1_IO_017 = tx_pin[1195];
  assign mb1_FA1_BB1_IO_016_mb1_FA2_BB1_IO_014 = tx_pin[1196];
  assign mb1_FA1_BB1_IO_017_mb1_FA2_BB1_IO_015 = tx_pin[1197];
  assign mb1_FA1_BB1_IO_018_mb1_FA2_BB1_IO_032 = tx_pin[1198];
  assign mb1_FA1_BB1_IO_019_mb1_FA2_BB1_IO_033 = tx_pin[1199];
  assign mb1_FA1_BB1_IO_020_mb1_FA2_BB1_IO_030 = tx_pin[1200];
  assign mb1_FA1_BB1_IO_021_mb1_FA2_BB1_IO_031 = tx_pin[1201];
  assign mb1_FA1_BB1_IO_022_mb1_FA2_BB1_IO_008 = tx_pin[1202];
  assign mb1_FA1_BB1_IO_023_mb1_FA2_BB1_IO_009 = tx_pin[1203];
  assign mb1_FA1_BB1_IO_024_mb1_FA2_BB1_IO_026 = tx_pin[1204];
  assign mb1_FA1_BB1_IO_025_mb1_FA2_BB1_IO_027 = tx_pin[1205];
  assign mb1_FA1_BB1_IO_026_mb1_FA2_BB1_IO_024 = tx_pin[1206];
  assign mb1_FA1_BB1_IO_027_mb1_FA2_BB1_IO_025 = tx_pin[1207];
  assign mb1_FA1_BB1_IO_028_mb1_FA2_BB1_IO_042 = tx_pin[1208];
  assign mb1_FA1_BB1_IO_029_mb1_FA2_BB1_IO_043 = tx_pin[1209];
  assign mb1_FA1_BB1_IO_030_mb1_FA2_BB1_IO_020 = tx_pin[1210];
  assign mb1_FA1_BB1_IO_031_mb1_FA2_BB1_IO_021 = tx_pin[1211];
  assign mb1_FA1_BB1_IO_032_mb1_FA2_BB1_IO_018 = tx_pin[1212];
  assign mb1_FA1_BB1_IO_033_mb1_FA2_BB1_IO_019 = tx_pin[1213];
  assign mb1_FA1_BB1_IO_034_mb1_FA2_BB1_IO_036 = tx_pin[1214];
  assign mb1_FA1_BB1_IO_035_mb1_FA2_BB1_IO_037 = tx_pin[1215];
  assign mb1_FA1_BB1_IO_036_mb1_FA2_BB1_IO_034 = tx_pin[1216];
  assign mb1_FA1_BB1_IO_037_mb1_FA2_BB1_IO_035 = tx_pin[1217];
  assign mb1_FA1_BB1_IO_038_mb1_FA2_BB1_IO_052 = tx_pin[1218];
  assign mb1_FA1_BB1_IO_039_mb1_FA2_BB1_IO_053 = tx_pin[1219];
  assign mb1_FA1_BB1_IO_040_mb1_FA2_BB1_IO_050 = tx_pin[1220];
  assign mb1_FA1_BB1_IO_041_mb1_FA2_BB1_IO_051 = tx_pin[1221];
  assign mb1_FA1_BB1_IO_042_mb1_FA2_BB1_IO_028 = tx_pin[1222];
  assign mb1_FA1_BB1_IO_043_mb1_FA2_BB1_IO_029 = tx_pin[1223];
  assign mb1_FA1_BB1_IO_044_mb1_FA2_BB1_IO_046 = tx_pin[1224];
  assign mb1_FA1_BB1_IO_045_mb1_FA2_BB1_IO_047 = tx_pin[1225];
  assign mb1_FA1_BB1_IO_046_mb1_FA2_BB1_IO_044 = tx_pin[1226];
  assign mb1_FA1_BB1_IO_047_mb1_FA2_BB1_IO_045 = tx_pin[1227];
  assign mb1_FA1_BB1_IO_048_mb1_FA2_BB1_IO_062 = tx_pin[1228];
  assign mb1_FA1_BB1_IO_049_mb1_FA2_BB1_IO_063 = tx_pin[1229];
  assign mb1_FA1_BB1_IO_050_mb1_FA2_BB1_IO_040 = tx_pin[1230];
  assign mb1_FA1_BB1_IO_051_mb1_FA2_BB1_IO_041 = tx_pin[1231];
  assign mb1_FA1_BB1_IO_052_mb1_FA2_BB1_IO_038 = tx_pin[1232];
  assign mb1_FA1_BB1_IO_053_mb1_FA2_BB1_IO_039 = tx_pin[1233];
  assign mb1_FA1_BB1_IO_054_mb1_FA2_BB1_IO_056 = tx_pin[1234];
  assign mb1_FA1_BB1_IO_055_mb1_FA2_BB1_IO_057 = tx_pin[1235];
  assign mb1_FA1_BB1_IO_056_mb1_FA2_BB1_IO_054 = tx_pin[1236];
  assign mb1_FA1_BB1_IO_057_mb1_FA2_BB1_IO_055 = tx_pin[1237];
  assign mb1_FA1_BB1_IO_058_mb1_FA2_BB1_IO_072 = tx_pin[1238];
  assign mb1_FA1_BB1_IO_059_mb1_FA2_BB1_IO_073 = tx_pin[1239];
  assign mb1_FA1_BB1_IO_060_mb1_FA2_BB1_IO_070 = tx_pin[1240];
  assign mb1_FA1_BB1_IO_061_mb1_FA2_BB1_IO_071 = tx_pin[1241];
  assign mb1_FA1_BB1_IO_062_mb1_FA2_BB1_IO_048 = tx_pin[1242];
  assign mb1_FA1_BB1_IO_063_mb1_FA2_BB1_IO_049 = tx_pin[1243];
  assign mb1_FA1_BB1_IO_064_mb1_FA2_BB1_IO_066 = tx_pin[1244];
  assign mb1_FA1_BB1_IO_065_mb1_FA2_BB1_IO_067 = tx_pin[1245];
  assign mb1_FA1_BB1_IO_066_mb1_FA2_BB1_IO_064 = tx_pin[1246];
  assign mb1_FA1_BB1_IO_067_mb1_FA2_BB1_IO_065 = tx_pin[1247];
  assign mb1_FA1_BB1_IO_068_mb1_FA2_BB1_IO_082 = tx_pin[1248];
  assign mb1_FA1_BB1_IO_069_mb1_FA2_BB1_IO_083 = tx_pin[1249];
  assign mb1_FA1_BB1_IO_070_mb1_FA2_BB1_IO_060 = tx_pin[1250];
  assign mb1_FA1_BB1_IO_071_mb1_FA2_BB1_IO_061 = tx_pin[1251];
  assign mb1_FA1_BB1_IO_072_mb1_FA2_BB1_IO_058 = tx_pin[1252];
  assign mb1_FA1_BB1_IO_073_mb1_FA2_BB1_IO_059 = tx_pin[1253];
  assign mb1_FA1_BB1_IO_074_mb1_FA2_BB1_IO_076 = tx_pin[1254];
  assign mb1_FA1_BB1_IO_075_mb1_FA2_BB1_IO_077 = tx_pin[1255];
  assign mb1_FA1_BB1_IO_076_mb1_FA2_BB1_IO_074 = tx_pin[1256];
  assign mb1_FA1_BB1_IO_077_mb1_FA2_BB1_IO_075 = tx_pin[1257];
  assign mb1_FA1_BB1_IO_078_mb1_FA2_BB1_IO_092 = tx_pin[1258];
  assign mb1_FA1_BB1_IO_079_mb1_FA2_BB1_IO_093 = tx_pin[1259];
  assign mb1_FA1_BB1_IO_080_mb1_FA2_BB1_IO_090 = tx_pin[1260];
  assign mb1_FA1_BB1_IO_081_mb1_FA2_BB1_IO_091 = tx_pin[1261];
  assign mb1_FA1_BB1_IO_082_mb1_FA2_BB1_IO_068 = tx_pin[1262];
  assign mb1_FA1_BB1_IO_083_mb1_FA2_BB1_IO_069 = tx_pin[1263];
  assign mb1_FA1_BB1_IO_084_mb1_FA2_BB1_IO_086 = tx_pin[1264];
  assign mb1_FA1_BB1_IO_085_mb1_FA2_BB1_IO_087 = tx_pin[1265];
  assign mb1_FA1_BB1_IO_086_mb1_FA2_BB1_IO_084 = tx_pin[1266];
  assign mb1_FA1_BB1_IO_087_mb1_FA2_BB1_IO_085 = tx_pin[1267];
  assign mb1_FA1_BB1_IO_088_mb1_FA2_BB1_IO_102 = tx_pin[1268];
  assign mb1_FA1_BB1_IO_089_mb1_FA2_BB1_IO_103 = tx_pin[1269];
  assign mb1_FA1_BB1_IO_090_mb1_FA2_BB1_IO_080 = tx_pin[1270];
  assign mb1_FA1_BB1_IO_091_mb1_FA2_BB1_IO_081 = tx_pin[1271];
  assign mb1_FA1_BB1_IO_092_mb1_FA2_BB1_IO_078 = tx_pin[1272];
  assign mb1_FA1_BB1_IO_093_mb1_FA2_BB1_IO_079 = tx_pin[1273];
  assign mb1_FA1_BB1_IO_094_mb1_FA2_BB1_IO_096 = tx_pin[1274];
  assign mb1_FA1_BB1_IO_095_mb1_FA2_BB1_IO_097 = tx_pin[1275];
  assign mb1_FA1_BB1_IO_096_mb1_FA2_BB1_IO_094 = tx_pin[1276];
  assign mb1_FA1_BB1_IO_097_mb1_FA2_BB1_IO_095 = tx_pin[1277];
  assign mb1_FA1_BB1_IO_098_mb1_FA2_BB1_IO_112 = tx_pin[1278];
  assign mb1_FA1_BB1_IO_099_mb1_FA2_BB1_IO_113 = tx_pin[1279];
  assign mb1_FA1_BB1_IO_100_mb1_FA2_BB1_IO_110 = tx_pin[1280];
  assign mb1_FA1_BB1_IO_101_mb1_FA2_BB1_IO_111 = tx_pin[1281];
  assign mb1_FA1_BB1_IO_102_mb1_FA2_BB1_IO_088 = tx_pin[1282];
  assign mb1_FA1_BB1_IO_103_mb1_FA2_BB1_IO_089 = tx_pin[1283];
  assign mb1_FA1_BB1_IO_104_mb1_FA2_BB1_IO_106 = tx_pin[1284];
  assign mb1_FA1_BB1_IO_105_mb1_FA2_BB1_IO_107 = tx_pin[1285];
  assign mb1_FA1_BB1_IO_106_mb1_FA2_BB1_IO_104 = tx_pin[1286];
  assign mb1_FA1_BB1_IO_107_mb1_FA2_BB1_IO_105 = tx_pin[1287];
  assign mb1_FA1_BB1_IO_108_mb1_FA2_BB1_IO_122 = tx_pin[1288];
  assign mb1_FA1_BB1_IO_109_mb1_FA2_BB1_IO_123 = tx_pin[1289];
  assign mb1_FA1_BB1_IO_110_mb1_FA2_BB1_IO_100 = tx_pin[1290];
  assign mb1_FA1_BB1_IO_111_mb1_FA2_BB1_IO_101 = tx_pin[1291];
  assign mb1_FA1_BB1_IO_112_mb1_FA2_BB1_IO_098 = tx_pin[1292];
  assign mb1_FA1_BB1_IO_113_mb1_FA2_BB1_IO_099 = tx_pin[1293];
  assign mb1_FA1_BB1_IO_114_mb1_FA2_BB1_IO_116 = tx_pin[1294];
  assign mb1_FA1_BB1_IO_115_mb1_FA2_BB1_IO_117 = tx_pin[1295];
  assign mb1_FA1_BB1_IO_116_mb1_FA2_BB1_IO_114 = tx_pin[1296];
  assign mb1_FA1_BB1_IO_117_mb1_FA2_BB1_IO_115 = tx_pin[1297];
  assign mb1_FA1_BB1_IO_118_mb1_FA2_BB1_IO_132 = tx_pin[1298];
  assign mb1_FA1_BB1_IO_119_mb1_FA2_BB1_IO_133 = tx_pin[1299];
  assign mb1_FA1_BB1_IO_120_mb1_FA2_BB1_IO_130 = tx_pin[1300];
  assign mb1_FA1_BB1_IO_121_mb1_FA2_BB1_IO_131 = tx_pin[1301];
  assign mb1_FA1_BB1_IO_122_mb1_FA2_BB1_IO_108 = tx_pin[1302];
  assign mb1_FA1_BB1_IO_123_mb1_FA2_BB1_IO_109 = tx_pin[1303];
  assign mb1_FA1_BB1_IO_124_mb1_FA2_BB1_IO_126 = tx_pin[1304];
  assign mb1_FA1_BB1_IO_125_mb1_FA2_BB1_IO_127 = tx_pin[1305];
  assign mb1_FA1_BB1_IO_126_mb1_FA2_BB1_IO_124 = tx_pin[1306];
  assign mb1_FA1_BB1_IO_127_mb1_FA2_BB1_IO_125 = tx_pin[1307];
  assign mb1_FA1_BB1_IO_130_mb1_FA2_BB1_IO_120 = tx_pin[1308];
  assign mb1_FA1_BB1_IO_131_mb1_FA2_BB1_IO_121 = tx_pin[1309];
  assign mb1_FA1_BB1_IO_132_mb1_FA2_BB1_IO_118 = tx_pin[1310];
  assign mb1_FA1_BB1_IO_133_mb1_FA2_BB1_IO_119 = tx_pin[1311];
  assign mb1_FA1_BB1_IO_134_mb1_FA2_BB1_IO_136 = tx_pin[1312];
  assign mb1_FA1_BB1_IO_136_mb1_FA2_BB1_IO_134 = tx_pin[1313];

  dbst # (
    .DEVICE             ( "XVUP"   ),
    .TX_PINS            ( TX_PINS               ),
    .RX_PINS            ( RX_PINS               ),
    .DIFF_ENABLED       ( 0 ),
    .USE_CLK_INPUT_BUFG ( USE_CLK_INPUT_BUFG    )
  ) U_DBST (
    .tx_pin        ( tx_pin      ),
    .tx_pin_p      (             ),
    .tx_pin_n      (             ),
    .rx_pin        ( '0          ),
    .rx_pin_p      ( '0          ),
    .rx_pin_n      ( '0          ),
    .clk_p         ( CLK_P[1:0]  ),
    .clk_n         ( CLK_N[1:0]  ),
    .sync_p        ( SYNC_P[1:0] ),
    .sync_n        ( SYNC_N[1:0] ),
    .dmbi_f2h_o    ( DMBI_F2H    ),
    .dmbi_h2f_i    ( DMBI_H2F    )
  );
  
endmodule
